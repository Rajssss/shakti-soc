/*
Copyright (c) 2019, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.
* Redistributions in binary form must reproduce the above copyright notice, this list of
  conditions and the following disclaimer in the documentation and/or other materials provided
 with the distribution.
* Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------
*/

/*
   This BSV file has been generated by the PinMux tool available at:
   https://bitbucket.org/casl/pinmux.

   Authors: Neel Gala, Luke
   Date of generation: Tue Jul  9 13:39:32 2019
*/

package pinmux;

  import GetPut::*;
  import Vector::*;

      (*always_ready,always_enabled*)
      interface MuxSelectionLines;

      // declare the method which will capture the user pin-mux
      // selection values.The width of the input is dependent on the number
      // of muxes happening per IO. For now we have a generalized width
      // where each IO will have the same number of muxes.
     method  Action cell7_mux (Bit#(2) in);
     method  Action cell8_mux (Bit#(2) in);
     method  Action cell9_mux (Bit#(2) in);
     method  Action cell10_mux (Bit#(2) in);
     method  Action cell12_mux (Bit#(2) in);
     method  Action cell13_mux (Bit#(2) in);
     method  Action cell16_mux (Bit#(2) in);
     method  Action cell17_mux (Bit#(2) in);
     method  Action cell18_mux (Bit#(2) in);
     method  Action cell19_mux (Bit#(2) in);
     method  Action cell20_mux (Bit#(2) in);
      endinterface


      interface IOCellSide;
      // declare the interface to the IO cells.
      // Each IO cell will have 1 input field (output from pin mux)
      // and an output and out-enable field (input to pinmux)
          // interface declaration between IO-7 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io7_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io7_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io7_cell_in (Bit#(1) in);
          // interface declaration between IO-8 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io8_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io8_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io8_cell_in (Bit#(1) in);
          // interface declaration between IO-9 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io9_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io9_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io9_cell_in (Bit#(1) in);
          // interface declaration between IO-10 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io10_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io10_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io10_cell_in (Bit#(1) in);
          // interface declaration between IO-12 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io12_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io12_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io12_cell_in (Bit#(1) in);
          // interface declaration between IO-13 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io13_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io13_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io13_cell_in (Bit#(1) in);
          // interface declaration between IO-16 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io16_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io16_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io16_cell_in (Bit#(1) in);
          // interface declaration between IO-17 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io17_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io17_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io17_cell_in (Bit#(1) in);
          // interface declaration between IO-18 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io18_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io18_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io18_cell_in (Bit#(1) in);
          // interface declaration between IO-19 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io19_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io19_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io19_cell_in (Bit#(1) in);
          // interface declaration between IO-20 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) io20_cell_out;
    (*always_ready,always_enabled*) method  Bit#(1) io20_cell_outen;
    (*always_ready,always_enabled,result="io"*) method
                       Action io20_cell_in (Bit#(1) in);
      endinterface

      // interface declaration between UART and pinmux
      (*always_ready,always_enabled*)
      interface PeripheralSideUART;
          interface Put#(Bit#(1)) tx;
          interface Get#(Bit#(1)) rx;
      endinterface

      // interface declaration between MSPI and pinmux
      (*always_ready,always_enabled*)
      interface PeripheralSideMSPI;
          interface Put#(Bit#(1)) clk;
          interface Put#(Bit#(1)) nss;
          interface Put#(Bit#(1)) mosi;
          interface Get#(Bit#(1)) miso;

      endinterface

      // interface declaration between GPIOA and pinmux
      (*always_ready,always_enabled*)
      interface PeripheralSideGPIOA;

          //interface Put#(Vector#(11,Bit#(1))) out;
          //interface Put#(Vector#(11,Bit#(1))) out_en;
          //interface Get#(Vector#(11,Bit#(1))) in;
          interface Put#(Bit#(11)) out;
          interface Put#(Bit#(11)) out_en;
          interface Get#(Bit#(11)) in;

      endinterface

      // interface declaration between PWM and pinmux
      (*always_ready,always_enabled*)
      interface PeripheralSidePWM;
          interface Put#(Bit#(1)) out;
      endinterface

      (*always_ready,always_enabled*)
      interface PeripheralSide;
      // declare the interface to the peripherals
      // Each peripheral's function will be either an input, output
      // or be bi-directional.  an input field will be an output from the
      // peripheral and an output field will be an input to the peripheral.
      // Bi-directional functions also have an output-enable (which
      // again comes *in* from the peripheral)
            interface PeripheralSideUART uart1;
            interface PeripheralSideUART uart2;
            interface PeripheralSideMSPI mspi;
            interface PeripheralSideGPIOA gpioa;
            interface PeripheralSidePWM pwm0;
            interface PeripheralSidePWM pwm1;
            interface PeripheralSidePWM pwm2;
            interface PeripheralSidePWM pwm3;
            interface PeripheralSidePWM pwm4;
            interface PeripheralSidePWM pwm5;
      endinterface


   interface Ifc_pinmux;
      // this interface controls how each IO cell is routed.  setting
      // any given IO cell's mux control value will result in redirection
      // of not just the input or output to different peripheral functions
      // but also the *direction* control - if appropriate - as well.
      interface MuxSelectionLines mux_lines;

      // this interface contains the inputs, outputs and direction-control
      // lines for all peripherals.  GPIO is considered to also be just
      // a peripheral because it also has in, out and direction-control.
      interface PeripheralSide peripheral_side;

      // this interface is to be linked to the individual IO cells.
      // if looking at a "non-muxed" GPIO design, basically the
      // IO cell input, output and direction-control wires are cut
      // (giving six pairs of dangling wires, named left and right)
      // these iocells are routed in their place on one side ("left")
      // and the matching *GPIO* peripheral interfaces in/out/dir
      // connect to the OTHER side ("right").  the result is that
      // the muxer settings end up controlling the routing of where
      // the I/O from the IOcell actually goes.
      interface IOCellSide iocell_side;
   endinterface

   (*synthesize*)
   module mkpinmux(Ifc_pinmux);

      // the followins wires capture the pin-mux selection
      // values for each mux assigned to a CELL

      Wire#(Bit#(2)) wrcell7_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell8_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell9_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell10_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell12_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell13_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell16_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell17_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell18_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell19_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell20_mux<-mkDWire(0);
      // following wires capture signals to IO CELL if io-7 is
      // allotted to it
      Wire#(Bit#(1)) cell7_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell7_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell7_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-8 is
      // allotted to it
      Wire#(Bit#(1)) cell8_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell8_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell8_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-9 is
      // allotted to it
      Wire#(Bit#(1)) cell9_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell9_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell9_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-10 is
      // allotted to it
      Wire#(Bit#(1)) cell10_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell10_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell10_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-12 is
      // allotted to it
      Wire#(Bit#(1)) cell12_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell12_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell12_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-13 is
      // allotted to it
      Wire#(Bit#(1)) cell13_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell13_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell13_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-16 is
      // allotted to it
      Wire#(Bit#(1)) cell16_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell16_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell16_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-17 is
      // allotted to it
      Wire#(Bit#(1)) cell17_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell17_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell17_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-18 is
      // allotted to it
      Wire#(Bit#(1)) cell18_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell18_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell18_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-19 is
      // allotted to it
      Wire#(Bit#(1)) cell19_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell19_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell19_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-20 is
      // allotted to it
      Wire#(Bit#(1)) cell20_mux_out<-mkDWire(0);
      Wire#(Bit#(1)) cell20_mux_outen<-mkDWire(0);
      Wire#(Bit#(1)) cell20_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if uart-1 is
      // allotted to it
      Wire#(Bit#(1)) wruart1_tx<-mkDWire(0);
      Wire#(Bit#(1)) wruart1_rx<-mkDWire(0);

      // following wires capture signals to IO CELL if uart-2 is
      // allotted to it
      Wire#(Bit#(1)) wruart2_tx<-mkDWire(0);
      Wire#(Bit#(1)) wruart2_rx<-mkDWire(0);

      // following wires capture signals to IO CELL if mspi-1 is
      // allotted to it
      Wire#(Bit#(1)) wrmspi2_clk<-mkDWire(0);
      Wire#(Bit#(1)) wrmspi2_nss<-mkDWire(0);
      Wire#(Bit#(1)) wrmspi2_mosi<-mkDWire(0);
      Wire#(Bit#(1)) wrmspi2_miso<-mkDWire(0);

      // following wires capture signals to IO CELL if gpioa-0 is
      // allotted to it
      Wire#(Bit#(1)) wrgpioa_a0_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a0_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a0_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a1_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a1_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a1_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a2_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a2_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a2_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a3_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a3_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a3_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a5_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a5_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a5_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a6_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a6_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a6_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a9_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a9_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a9_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a10_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a10_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a10_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a11_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a11_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a11_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a12_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a12_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a12_in<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a13_out<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a13_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrgpioa_a13_in<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-0 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm0_out<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-1 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm1_out<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-2 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm2_out<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-3 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm3_out<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-4 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm4_out<-mkDWire(0);

      // following wires capture signals to IO CELL if pwm-5 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm5_out<-mkDWire(0);


      /*====== This where the muxing starts for each io-cell======*/
      Wire#(Bit#(1)) val0<-mkDWire(0); // need a zero
      Wire#(Bit#(1)) val1<-mkDWire(1); // need a one
       // --------------------
      // ----- cell 7 -----

      // output muxer for cell idx 7
      cell7_mux_out=
			wrcell7_mux==0?wrgpioa_a0_out:
			wrcell7_mux==1?val0:
			wrcell7_mux==2?val0: // unused
			val0; // unused

      // outen muxer for cell idx 7
      cell7_mux_outen=
			wrcell7_mux==0?wrgpioa_a0_outen: // bi-directional
			wrcell7_mux==1?val1: // uart1_rx is an input
			wrcell7_mux==2?val0: // unused
			val0; // unused

      // priority-in-muxer for cell idx 0
      rule assign_wrgpioa_a0_in_on_cell7(wrcell7_mux==0);
        wrgpioa_a0_in<=cell7_mux_in;
        wruart1_rx<=val1;
      endrule

      rule assign_wruart1_rx_on_cell7(wrcell7_mux==1);
        wruart1_rx<=cell7_mux_in;
        wrgpioa_a0_in<=val0;
      endrule

      rule assign_wr_on_cell7_2(wrcell7_mux==2);
        wruart1_rx<=val1;
        wrgpioa_a0_in<=val0;
      endrule

      rule assign_wr_on_cell7_3(wrcell7_mux==3);
        wruart1_rx<=val1;
        wrgpioa_a0_in<=val0;
      endrule

      // --------------------
      // ----- cell 8 -----

      // output muxer for cell idx 8
      cell8_mux_out=
			wrcell8_mux==0?wrgpioa_a1_out:
			wrcell8_mux==1?wruart1_tx: // uart1_tx is an output
			wrcell8_mux==2?val0: // unused
			val0; // unused

      // outen muxer for cell idx 1
      cell8_mux_outen=
			wrcell8_mux==0?wrgpioa_a1_outen: // bi-directional
			wrcell8_mux==1?val0: // uart1_tx is an output
			wrcell8_mux==2?val0: // unused
			val0; // unused

      // priority-in-muxer for cell idx 8
      rule assign_wrgpioa_a1_in_on_cell8(wrcell8_mux==0);
        wrgpioa_a1_in<=cell8_mux_in;
      endrule

      rule assign_wr_on_cell8_1(wrcell8_mux==1);
        wrgpioa_a1_in<=val0;
      endrule

      rule assign_wr_on_cell8_2(wrcell8_mux==2);
        wrgpioa_a1_in<=val0;
      endrule

      rule assign_wr_on_cell8_3(wrcell8_mux==3);
        wrgpioa_a1_in<=val0;
      endrule

      // --------------------
      // ----- cell 9 -----

      // output muxer for cell idx 9
      cell9_mux_out=
			wrcell9_mux==0?wrgpioa_a2_out:
			wrcell9_mux==1?val0:
			wrcell9_mux==2?val0:
			val0; // unused

      // outen muxer for cell idx 9
      cell9_mux_outen=
			wrcell9_mux==0?wrgpioa_a2_outen: // bi-directional
			wrcell9_mux==1?val1: // uart2_rx is an input
			wrcell9_mux==2?val0:
			val0; // unused

      // priority-in-muxer for cell idx 2
      rule assign_wrgpioa_a2_in_on_cell9(wrcell9_mux==0);
        wrgpioa_a2_in<=cell9_mux_in;
        wruart2_rx<=val1;
      endrule

      rule assign_wruart2_rx_on_cell9(wrcell9_mux==1);
        wrgpioa_a2_in<=val0;
        wruart2_rx<=cell9_mux_in;
      endrule

      rule assign_wr_on_cell9_2(wrcell9_mux==2);
        wrgpioa_a2_in<=val0;
        wruart2_rx<=val1;
      endrule

      rule assign_wr_on_cell9_3(wrcell9_mux==3);
        wrgpioa_a2_in<=val0;
        wruart2_rx<=val1;
      endrule

      // --------------------
      // ----- cell 10 -----

      // output muxer for cell idx 10
      cell10_mux_out=
			wrcell10_mux==0?wrgpioa_a3_out:
			wrcell10_mux==1?wruart2_tx: // uart2_tx is an output
			wrcell10_mux==2?wrpwm0_out: // pwm0 is a output
			val0; // unused

      // outen muxer for cell idx 3
      cell10_mux_outen=
			wrcell10_mux==0?wrgpioa_a3_outen: // bi-directional
			wrcell10_mux==1?val0: // uart2_tx is an output
			wrcell10_mux==2?val0: // pwm0 is a output
			val0; // unused

      // priority-in-muxer for cell idx 3
      rule assign_wrgpioa_a3_in_on_cell10(wrcell10_mux==0);
        wrgpioa_a3_in<=cell10_mux_in;
      endrule

      rule assign_wr_on_cell10_1(wrcell10_mux==1);
        wrgpioa_a3_in<=val0;
      endrule

      rule assign_wr_on_cell10_2(wrcell10_mux==2);
        wrgpioa_a3_in<=val0;
      endrule

      rule assign_wr_on_cell10_3(wrcell10_mux==3);
        wrgpioa_a3_in<=val0;
      endrule

      // --------------------
      // --------------------
      // ----- cell 12 -----

      // output muxer for cell idx 12
      cell12_mux_out=
			wrcell12_mux==0?wrgpioa_a5_out:
			wrcell12_mux==1?val0: // unused
			wrcell12_mux==2?wrpwm1_out:
			val0; // unused

      // outen muxer for cell idx 12
      cell12_mux_outen=
			wrcell12_mux==0?wrgpioa_a5_outen: // bi-directional
			wrcell12_mux==1?val0: // unused
			wrcell12_mux==2?val0: // pwm1_out is an output
			val0; // unused

      // priority-in-muxer for cell idx 4
      rule assign_wrgpioa_a5_in_on_cell12(wrcell12_mux==0);
        wrgpioa_a5_in<=cell12_mux_in;
      endrule

      rule assign_wr_on_cell12_1(wrcell12_mux==1);
        wrgpioa_a5_in<=val0;
      endrule

      rule assign_wr_on_cell12_2(wrcell12_mux==2);
        wrgpioa_a5_in<=val0;
      endrule

      rule assign_wr_on_cell12_3(wrcell12_mux==3);
        wrgpioa_a5_in<=val0;
      endrule

      // --------------------
      // ----- cell 13 -----

      // output muxer for cell idx 13
      cell13_mux_out=
			wrcell13_mux==0?wrgpioa_a6_out:
			wrcell13_mux==1?val0: // unused
			wrcell13_mux==2?wrpwm2_out: // pwm2_out is an output
			val0; // unused

      // outen muxer for cell idx 13
      cell13_mux_outen=
			wrcell13_mux==0?wrgpioa_a6_outen: // bi-directional
			wrcell13_mux==1?val0: // unused
			wrcell13_mux==2?val0: // pwm2_out is an output
			val0; // unused

      // priority-in-muxer for cell idx 13
      rule assign_wrgpioa_a6_in_on_cell13(wrcell13_mux==0);
        wrgpioa_a6_in<=cell13_mux_in;
      endrule

      rule assign_wr_on_cell13_1(wrcell13_mux==1);
        wrgpioa_a6_in<=val0;
      endrule

      rule assign_wr_on_cell13_2(wrcell13_mux==2);
        wrgpioa_a6_in<=val0;
      endrule

      rule assign_wr_on_cell13_3(wrcell13_mux==3);
        wrgpioa_a6_in<=val0;
      endrule

      // --------------------
      // ----- cell 16 -----

      // output muxer for cell idx 16
      cell16_mux_out=
			wrcell16_mux==0?wrgpioa_a9_out:
			wrcell16_mux==1?val0: // unused
			wrcell16_mux==2?wrpwm3_out: // pwm3_out is an output
			val0; // unused

      // outen muxer for cell idx 16
      cell16_mux_outen=
			wrcell16_mux==0?wrgpioa_a9_outen: // bi-directional
			wrcell16_mux==1?val0: // unused
			wrcell16_mux==2?val0: // pwm3_out is an output
			val0; // unused

      // priority-in-muxer for cell idx 16
      rule assign_wrgpioa_a9_in_on_cell16(wrcell16_mux==0);
        wrgpioa_a9_in<=cell16_mux_in;
      endrule

      rule assign_wr_on_cell16_1(wrcell16_mux==1);
        wrgpioa_a9_in<=val0;
      endrule

      rule assign_wr_on_cell16_2(wrcell16_mux==2);
        wrgpioa_a9_in<=val0;
      endrule

      rule assign_wr_on_cell16_3(wrcell16_mux==3);
        wrgpioa_a9_in<=val0;
      endrule

      // --------------------
      // ----- cell 17 -----

      // output muxer for cell idx 17
      cell17_mux_out=
			wrcell17_mux==0?wrgpioa_a10_out:
			wrcell17_mux==1?wrmspi2_nss: // mspi nss is an output
			wrcell17_mux==2?wrpwm4_out: // pwm4_out is an output
			val0; // unused

      // outen muxer for cell idx 17
      cell17_mux_outen=
			wrcell17_mux==0?wrgpioa_a10_outen: // bi-directional
			wrcell17_mux==1?val0: // mspi_nss is an output
			wrcell17_mux==2?val0: // pwm4_out is an output
			val0; // unused

      // priority-in-muxer for cell idx 17
      rule assign_wrgpioa_a10_in_on_cell17(wrcell17_mux==0);
        wrgpioa_a10_in<=cell17_mux_in;
      endrule

      rule assign_wr_on_cell17_1(wrcell17_mux==1);
        wrgpioa_a10_in<=val0;
      endrule

      rule assign_wr_on_cell17_2(wrcell17_mux==2);
        wrgpioa_a10_in<=val0;
      endrule

      rule assign_wr_on_cell17_3(wrcell17_mux==3);
        wrgpioa_a10_in<=val0;
      endrule

      // --------------------
      // ----- cell 18 -----

      // output muxer for cell idx 18
      cell18_mux_out=
			wrcell18_mux==0?wrgpioa_a11_out:
			wrcell18_mux==1?wrmspi2_mosi:
			wrcell18_mux==2?wrpwm5_out:
			val0; // unused

      // outen muxer for cell idx 18
      cell18_mux_outen=
			wrcell18_mux==0?wrgpioa_a11_outen: // bi-directional
			wrcell18_mux==1?val0: // mspi1_mosi is an output
			wrcell18_mux==2?val0: // pwm4_out is an output
			val0; // unused

      // priority-in-muxer for cell idx 18
      rule assign_wrgpioa_a11_in_on_cell18(wrcell18_mux==0);
        wrgpioa_a11_in<=cell18_mux_in;
      endrule

      rule assign_wr_on_cell18_1(wrcell18_mux==1);
        wrgpioa_a11_in<=val0;
      endrule

      rule assign_wr_on_cell18_2(wrcell18_mux==2);
        wrgpioa_a11_in<=val0;
      endrule

      rule assign_wr_on_cell18_3(wrcell18_mux==3);
        wrgpioa_a11_in<=val0;
      endrule

      // --------------------
      // ----- cell 19 -----

      // output muxer for cell idx 19
      cell19_mux_out=
			wrcell19_mux==0?wrgpioa_a12_out:
			wrcell19_mux==1?val0: //mspi2_miso is an input
			wrcell19_mux==2?val0: // unused
			val0; // unused

      // outen muxer for cell idx 19
      cell19_mux_outen=
			wrcell19_mux==0?wrgpioa_a12_outen: // bi-directional
			wrcell19_mux==1?val1: // mspi2_miso is an input
			wrcell19_mux==2?val0: // unused
			val0; // unused

      // priority-in-muxer for cell idx 19
      rule assign_wrgpioa_a12_in_on_cell19(wrcell19_mux==0);
        wrgpioa_a12_in<=cell19_mux_in;
        wrmspi2_miso <=val0;
      endrule

      rule assign_wrmspi2_miso_in_on_cell19(wrcell19_mux==1);
        wrgpioa_a12_in<=val0;
        wrmspi2_miso <=cell19_mux_in;
      endrule

      rule assign_wr_on_cell19_2(wrcell19_mux==2);
        wrgpioa_a12_in<=val0;
        wrmspi2_miso <=val0;
      endrule

      rule assign_wr_on_cell19_3(wrcell19_mux==3);
        wrgpioa_a12_in<=val0;
        wrmspi2_miso <=val0;
      endrule

      // --------------------
      // ----- cell 20 -----

      // output muxer for cell idx 20
      cell20_mux_out=
			wrcell20_mux==0?wrgpioa_a13_out:
			wrcell20_mux==1?wrmspi2_clk: // mspi2_clk is an output
			wrcell20_mux==2?val0:
			val0; // unused

      // outen muxer for cell idx 20
      cell20_mux_outen=
			wrcell20_mux==0?wrgpioa_a13_outen: // bi-directional
			wrcell20_mux==1?val0: // dedicated output
			wrcell20_mux==2?val0:
			val0; // unused

      // priority-in-muxer for cell idx 20
      rule assign_wrgpioa_a13_in_on_cell20(wrcell20_mux==0);
        wrgpioa_a13_in<=cell20_mux_in;
      endrule

      rule assign_wr_on_cell20_1(wrcell20_mux==1);
        wrgpioa_a13_in<=val0;
      endrule

      rule assign_wr_on_cell20_2(wrcell20_mux==2);
        wrgpioa_a13_in<=val0;
      endrule

      rule assign_wr_on_cell20_3(wrcell20_mux==3);
        wrgpioa_a13_in<=val0;
      endrule

      /*=========================================*/
      // dedicated cells


      /*============================================================*/

  //interface pinmux_io = interface Ifc_pinmux

    interface mux_lines = interface MuxSelectionLines

      method Action  cell7_mux(Bit#(2) in);
         wrcell7_mux<=in;
      endmethod

      method Action  cell8_mux(Bit#(2) in);
         wrcell8_mux<=in;
      endmethod

      method Action  cell9_mux(Bit#(2) in);
         wrcell9_mux<=in;
      endmethod

      method Action  cell10_mux(Bit#(2) in);
         wrcell10_mux<=in;
      endmethod

      method Action  cell12_mux(Bit#(2) in);
         wrcell12_mux<=in;
      endmethod

      method Action  cell13_mux(Bit#(2) in);
         wrcell13_mux<=in;
      endmethod

      method Action  cell16_mux(Bit#(2) in);
         wrcell16_mux<=in;
      endmethod

      method Action  cell17_mux(Bit#(2) in);
         wrcell17_mux<=in;
      endmethod

      method Action  cell18_mux(Bit#(2) in);
         wrcell18_mux<=in;
      endmethod

      method Action  cell19_mux(Bit#(2) in);
         wrcell19_mux<=in;
      endmethod

      method Action  cell20_mux(Bit#(2) in);
         wrcell20_mux<=in;
      endmethod

    endinterface;

    interface iocell_side = interface IOCellSide

      method io7_cell_out=cell7_mux_out;
      method io7_cell_outen=cell7_mux_outen;
      method Action  io7_cell_in(Bit#(1) in);
         cell7_mux_in<=in;
      endmethod

      method io8_cell_out=cell8_mux_out;
      method io8_cell_outen=cell8_mux_outen;
      method Action  io8_cell_in(Bit#(1) in);
         cell8_mux_in<=in;
      endmethod

      method io9_cell_out=cell9_mux_out;
      method io9_cell_outen=cell9_mux_outen;
      method Action  io9_cell_in(Bit#(1) in);
         cell9_mux_in<=in;
      endmethod

      method io10_cell_out=cell10_mux_out;
      method io10_cell_outen=cell10_mux_outen;
      method Action  io10_cell_in(Bit#(1) in);
         cell10_mux_in<=in;
      endmethod

      method io12_cell_out=cell12_mux_out;
      method io12_cell_outen=cell12_mux_outen;
      method Action  io12_cell_in(Bit#(1) in);
         cell12_mux_in<=in;
      endmethod

      method io13_cell_out=cell13_mux_out;
      method io13_cell_outen=cell13_mux_outen;
      method Action  io13_cell_in(Bit#(1) in);
         cell13_mux_in<=in;
      endmethod

      method io16_cell_out=cell16_mux_out;
      method io16_cell_outen=cell16_mux_outen;
      method Action  io16_cell_in(Bit#(1) in);
         cell16_mux_in<=in;
      endmethod

      method io17_cell_out=cell17_mux_out;
      method io17_cell_outen=cell17_mux_outen;
      method Action  io17_cell_in(Bit#(1) in);
         cell17_mux_in<=in;
      endmethod

      method io18_cell_out=cell18_mux_out;
      method io18_cell_outen=cell18_mux_outen;
      method Action  io18_cell_in(Bit#(1) in);
         cell18_mux_in<=in;
      endmethod

      method io19_cell_out=cell19_mux_out;
      method io19_cell_outen=cell19_mux_outen;
      method Action  io19_cell_in(Bit#(1) in);
         cell19_mux_in<=in;
      endmethod

      method io20_cell_out=cell20_mux_out;
      method io20_cell_outen=cell20_mux_outen;
      method Action  io20_cell_in(Bit#(1) in);
         cell20_mux_in<=in;
      endmethod

     endinterface;

     interface peripheral_side = interface PeripheralSide
        interface uart1 = interface PeripheralSideUART
            interface tx = interface Put
              method Action put(Bit#(1) in);
                wruart1_tx<=in;
              endmethod
            endinterface;
            interface rx = interface Get
              method ActionValue#(Bit#(1)) get;
                return wruart1_rx;
              endmethod
            endinterface;
        endinterface;

        interface uart2 = interface PeripheralSideUART
            interface tx = interface Put
              method Action put(Bit#(1) in);
                wruart2_tx<=in;
              endmethod
            endinterface;
            interface rx = interface Get
              method ActionValue#(Bit#(1)) get;
                return wruart2_rx;
              endmethod
            endinterface;
        endinterface;

        interface mspi = interface PeripheralSideMSPI
            interface clk = interface Put
              method Action put(Bit#(1) in);
                wrmspi2_clk<=in;
              endmethod
            endinterface;
            interface nss = interface Put
              method Action put(Bit#(1) in);
                wrmspi2_nss<=in;
              endmethod
            endinterface;
              interface mosi = interface Put
                 method Action put(Bit#(1) in);
                   wrmspi2_mosi <= in;
                 endmethod
               endinterface;
               interface miso = interface Get
                 method ActionValue#(Bit#(1)) get;
                   Bit#(1) tget;
                   tget = wrmspi2_miso;
                   return tget;
                 endmethod
               endinterface;

        endinterface;

        interface gpioa = interface PeripheralSideGPIOA

              interface out = interface Put#(11)
                 //method Action put(Vector#(11,Bit#(1)) in);
                 method Action put(Bit#(11) in);
                   wrgpioa_a0_out <= in[0];
                   wrgpioa_a1_out <= in[1];
                   wrgpioa_a2_out <= in[2];
                   wrgpioa_a3_out <= in[3];
                   wrgpioa_a5_out <= in[4];
                   wrgpioa_a6_out <= in[5];
                   wrgpioa_a9_out <= in[6];
                   wrgpioa_a10_out <= in[7];
                   wrgpioa_a11_out <= in[8];
                   wrgpioa_a12_out <= in[9];
                   wrgpioa_a13_out <= in[10];
                 endmethod
               endinterface;
               interface out_en = interface Put#(11)
                 //method Action put(Vector#(11,Bit#(1)) in);
                 method Action put(Bit#(11) in);
                   wrgpioa_a0_outen <= ~in[0];
                   wrgpioa_a1_outen <= ~in[1];
                   wrgpioa_a2_outen <= ~in[2];
                   wrgpioa_a3_outen <= ~in[3];
                   wrgpioa_a5_outen <= ~in[4];
                   wrgpioa_a6_outen <= ~in[5];
                   wrgpioa_a9_outen <= ~in[6];
                   wrgpioa_a10_outen <= ~in[7];
                   wrgpioa_a11_outen <= ~in[8];
                   wrgpioa_a12_outen <= ~in[9];
                   wrgpioa_a13_outen <= ~in[10];
                 endmethod
               endinterface;
               interface in = interface Get#(11)
                 //method ActionValue#(Vector#(11,Bit#(1))) get;
                 method ActionValue#(Bit#(11)) get;
                   //Vector#(11,Bit#(1)) tget;
                   Bit#(11) tget;
                   tget[0] = wrgpioa_a0_in;
                   tget[1] = wrgpioa_a1_in;
                   tget[2] = wrgpioa_a2_in;
                   tget[3] = wrgpioa_a3_in;
                   tget[4] = wrgpioa_a5_in;
                   tget[5] = wrgpioa_a6_in;
                   tget[6] = wrgpioa_a9_in;
                   tget[7] = wrgpioa_a10_in;
                   tget[8] = wrgpioa_a11_in;
                   tget[9] = wrgpioa_a12_in;
                   tget[10] = wrgpioa_a13_in;
                   return tget;
                 endmethod
               endinterface;

        endinterface;

        interface pwm0 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm0_out<=in;
              endmethod
            endinterface;
        endinterface;

        interface pwm1 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm1_out<=in;
              endmethod
            endinterface;
        endinterface;

        interface pwm2 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm2_out<=in;
              endmethod
            endinterface;
        endinterface;

        interface pwm3 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm3_out<=in;
              endmethod
            endinterface;
        endinterface;

        interface pwm4 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm4_out<=in;
              endmethod
            endinterface;
        endinterface;

        interface pwm5 = interface PeripheralSidePWM
            interface out = interface Put
              method Action put(Bit#(1) in);
                wrpwm5_out<=in;
              endmethod
            endinterface;
        endinterface;


      endinterface;
   endmodule
endpackage
