// Bluespec wrapper, created by Import BVI Wizard
// Created on: Mon Dec 02 14:47:41 IST 2019
// Created by: shakti6
// Bluespec version: 2019.05.beta2 2019-05-24 a88bf40db


interface Ifc_aardonyx_wrapper;

  interface Inout#(Bit#(1)) gpio_0;
	interface Inout#(Bit(#1)) gpio_1;
	interface Inout#(Bit(#1)) gpio_2;
	interface Inout#(Bit(#1)) gpio_3;
	interface Inout#(Bit(#1)) gpio_4;
	interface Inout#(Bit(#1)) gpio_5;
	interface Inout#(Bit(#1)) gpio_6;
	interface Inout#(Bit(#1)) gpio_7;
	interface Inout#(Bit(#1)) gpio_8;
	interface Inout#(Bit(#1)) gpio_9;
	interface Inout#(Bit(#1)) gpio_10;
	interface Inout#(Bit(#1)) gpio_11;
	interface Inout#(Bit(#1)) gpio_12;
	interface Inout#(Bit(#1)) gpio_13;
	interface Inout#(Bit(#1)) gpio_14;
	interface Inout#(Bit(#1)) gpio_15;
	interface Inout#(Bit(#1)) i2c1_scl;
	interface Inout#(Bit(#1)) i2c1_sda;
	interface Inout#(Bit(#1)) qspi0_io0;
	interface Inout#(Bit(#1)) qspi0_io1;
	interface Inout#(Bit(#1)) qspi0_io2;
	interface Inout#(Bit(#1)) qspi0_io3;
	interface Inout#(Bit(#1)) i2c0_sda;
	interface Inout#(Bit(#1)) i2c0_scl;
	interface Inout#(Bit(#1)) sdram_d0;
	interface Inout#(Bit(#1)) sdram_d1;
	interface Inout#(Bit(#1)) sdram_d2;
	interface Inout#(Bit(#1)) sdram_d3;
	interface Inout#(Bit(#1)) sdram_d4;
	interface Inout#(Bit(#1)) sdram_d5;
	interface Inout#(Bit(#1)) sdram_d6;
	interface Inout#(Bit(#1)) sdram_d7;
	interface Inout#(Bit(#1)) sdram_d8;
	interface Inout#(Bit(#1)) sdram_d9;
	interface Inout#(Bit(#1)) sdram_d10;
	interface Inout#(Bit(#1)) sdram_d11;
	interface Inout#(Bit(#1)) sdram_d12;
	interface Inout#(Bit(#1)) sdram_d13;
	interface Inout#(Bit(#1)) sdram_d14;
	interface Inout#(Bit(#1)) sdram_d15;
	interface Inout#(Bit(#1)) sdram_d16;
	interface Inout#(Bit(#1)) sdram_d17;
	interface Inout#(Bit(#1)) sdram_d18;
	interface Inout#(Bit(#1)) sdram_d19;
	interface Inout#(Bit(#1)) sdram_d20;
	interface Inout#(Bit(#1)) sdram_d21;
	interface Inout#(Bit(#1)) sdram_d22;
	interface Inout#(Bit(#1)) sdram_d23;
	interface Inout#(Bit(#1)) sdram_d24;
	interface Inout#(Bit(#1)) sdram_d25;
	interface Inout#(Bit(#1)) sdram_d26;
	interface Inout#(Bit(#1)) sdram_d27;
	interface Inout#(Bit(#1)) sdram_d28;
	interface Inout#(Bit(#1)) sdram_d29;
	interface Inout#(Bit(#1)) sdram_d30;
	interface Inout#(Bit(#1)) sdram_d31;
	method Action ispi0_miso ();
	method Action iuart0_rx ();
	method Action itms ();
	method Action itrst ();
	method Action itck ();
	method Action itdi ();
	method Action ispi1_miso ();
	method Action iboot_mode0 ();
	method Action iboot_mode1 ();
	method Action itest_mode ();
	method Bool ospi0_ncs ();
	method Bool ospi0_clk ();
	method Bool ospi0_mosi ();
	method Bool oqspi0_clk ();
	method Bool oqspi0_ncs ();
	method Bool ouart0_tx ();
	method Bool otdo ();
	method Bool osdram_a0 ();
	method Bool osdram_a1 ();
	method Bool osdram_a2 ();
	method Bool osdram_a3 ();
	method Bool osdram_a4 ();
	method Bool osdram_a5 ();
	method Bool osdram_a6 ();
	method Bool osdram_a7 ();
	method Bool osdram_a8 ();
	method Bool osdram_a9 ();
	method Bool osdram_a10 ();
	method Bool osdram_a11 ();
	method Bool osdram_a12 ();
	method Bool osdram_dq0 ();
	method Bool osdram_dq1 ();
	method Bool osdram_dq2 ();
	method Bool osdram_dq3 ();
	method Bool osdram_ba0 ();
	method Bool osdram_ba1 ();
	method Bool osdram_cs ();
	method Bool osdram_ras ();
	method Bool osdram_cas ();
	method Bool osdram_we ();
	method Bool osdram_clk ();
	method Bool osdram_cke ();
	method Bool ospi1_ncs ();
	method Bool ospi1_clk ();
	method Bool ospi1_mosi ();
endinterface

import "BVI" aardonyx_wrapper =
module mkaardonyx_wrapper  (Ifc_aardonyx_wrapper);

	default_clock clk_clk;
	default_reset rst_reset;

	input_clock clk_clk (clk)  <- exposeCurrentClock;
	input_reset rst_reset (reset) clocked_by(clk_clk)  <- exposeCurrentReset;


	method ispi0_miso ()
		 enable(spi0_miso) clocked_by(clk_clk) reset_by(rst_reset);
	method iuart0_rx ()
		 enable(uart0_rx) clocked_by(clk_clk) reset_by(rst_reset);
	method itms ()
		 enable(tms) clocked_by(clk_clk) reset_by(rst_reset);
	method itrst ()
		 enable(trst) clocked_by(clk_clk) reset_by(rst_reset);
	method itck ()
		 enable(tck) clocked_by(clk_clk) reset_by(rst_reset);
	method itdi ()
		 enable(tdi) clocked_by(clk_clk) reset_by(rst_reset);
	method ispi1_miso ()
		 enable(spi1_miso) clocked_by(clk_clk) reset_by(rst_reset);
	method iboot_mode0 ()
		 enable(boot_mode0) clocked_by(clk_clk) reset_by(rst_reset);
	method iboot_mode1 ()
		 enable(boot_mode1) clocked_by(clk_clk) reset_by(rst_reset);
	method itest_mode ()
		 enable(test_mode) clocked_by(clk_clk) reset_by(rst_reset);
	method spi0_ncs ospi0_ncs ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method spi0_clk ospi0_clk ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method spi0_mosi ospi0_mosi ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method qspi0_clk oqspi0_clk ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method qspi0_ncs oqspi0_ncs ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method uart0_tx ouart0_tx ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method tdo otdo ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a0 osdram_a0 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a1 osdram_a1 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a2 osdram_a2 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a3 osdram_a3 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a4 osdram_a4 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a5 osdram_a5 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a6 osdram_a6 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a7 osdram_a7 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a8 osdram_a8 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a9 osdram_a9 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a10 osdram_a10 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a11 osdram_a11 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_a12 osdram_a12 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_dq0 osdram_dq0 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_dq1 osdram_dq1 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_dq2 osdram_dq2 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_dq3 osdram_dq3 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_ba0 osdram_ba0 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_ba1 osdram_ba1 ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_cs osdram_cs ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_ras osdram_ras ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_cas osdram_cas ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_we osdram_we ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_clk osdram_clk ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method sdram_cke osdram_cke ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method spi1_ncs ospi1_ncs ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method spi1_clk ospi1_clk ()
		 clocked_by(clk_clk) reset_by(rst_reset);
	method spi1_mosi ospi1_mosi ()
		 clocked_by(clk_clk) reset_by(rst_reset);

	schedule ispi0_miso C ispi0_miso;
	schedule ispi0_miso CF iuart0_rx;
	schedule ispi0_miso CF itms;
	schedule ispi0_miso CF itrst;
	schedule ispi0_miso CF itck;
	schedule ispi0_miso CF itdi;
	schedule ispi0_miso CF ispi1_miso;
	schedule ispi0_miso CF iboot_mode0;
	schedule ispi0_miso CF iboot_mode1;
	schedule ispi0_miso CF itest_mode;
	schedule ospi0_ncs SB ispi0_miso;
	schedule ospi0_clk SB ispi0_miso;
	schedule ospi0_mosi SB ispi0_miso;
	schedule oqspi0_clk SB ispi0_miso;
	schedule oqspi0_ncs SB ispi0_miso;
	schedule ouart0_tx SB ispi0_miso;
	schedule otdo SB ispi0_miso;
	schedule osdram_a0 SB ispi0_miso;
	schedule osdram_a1 SB ispi0_miso;
	schedule osdram_a2 SB ispi0_miso;
	schedule osdram_a3 SB ispi0_miso;
	schedule osdram_a4 SB ispi0_miso;
	schedule osdram_a5 SB ispi0_miso;
	schedule osdram_a6 SB ispi0_miso;
	schedule osdram_a7 SB ispi0_miso;
	schedule osdram_a8 SB ispi0_miso;
	schedule osdram_a9 SB ispi0_miso;
	schedule osdram_a10 SB ispi0_miso;
	schedule osdram_a11 SB ispi0_miso;
	schedule osdram_a12 SB ispi0_miso;
	schedule osdram_dq0 SB ispi0_miso;
	schedule osdram_dq1 SB ispi0_miso;
	schedule osdram_dq2 SB ispi0_miso;
	schedule osdram_dq3 SB ispi0_miso;
	schedule osdram_ba0 SB ispi0_miso;
	schedule osdram_ba1 SB ispi0_miso;
	schedule osdram_cs SB ispi0_miso;
	schedule osdram_ras SB ispi0_miso;
	schedule osdram_cas SB ispi0_miso;
	schedule osdram_we SB ispi0_miso;
	schedule osdram_clk SB ispi0_miso;
	schedule osdram_cke SB ispi0_miso;
	schedule ospi1_ncs SB ispi0_miso;
	schedule ospi1_clk SB ispi0_miso;
	schedule ospi1_mosi SB ispi0_miso;
	schedule iuart0_rx C iuart0_rx;
	schedule iuart0_rx CF itms;
	schedule iuart0_rx CF itrst;
	schedule iuart0_rx CF itck;
	schedule iuart0_rx CF itdi;
	schedule iuart0_rx CF ispi1_miso;
	schedule iuart0_rx CF iboot_mode0;
	schedule iuart0_rx CF iboot_mode1;
	schedule iuart0_rx CF itest_mode;
	schedule ospi0_ncs SB iuart0_rx;
	schedule ospi0_clk SB iuart0_rx;
	schedule ospi0_mosi SB iuart0_rx;
	schedule oqspi0_clk SB iuart0_rx;
	schedule oqspi0_ncs SB iuart0_rx;
	schedule ouart0_tx SB iuart0_rx;
	schedule otdo SB iuart0_rx;
	schedule osdram_a0 SB iuart0_rx;
	schedule osdram_a1 SB iuart0_rx;
	schedule osdram_a2 SB iuart0_rx;
	schedule osdram_a3 SB iuart0_rx;
	schedule osdram_a4 SB iuart0_rx;
	schedule osdram_a5 SB iuart0_rx;
	schedule osdram_a6 SB iuart0_rx;
	schedule osdram_a7 SB iuart0_rx;
	schedule osdram_a8 SB iuart0_rx;
	schedule osdram_a9 SB iuart0_rx;
	schedule osdram_a10 SB iuart0_rx;
	schedule osdram_a11 SB iuart0_rx;
	schedule osdram_a12 SB iuart0_rx;
	schedule osdram_dq0 SB iuart0_rx;
	schedule osdram_dq1 SB iuart0_rx;
	schedule osdram_dq2 SB iuart0_rx;
	schedule osdram_dq3 SB iuart0_rx;
	schedule osdram_ba0 SB iuart0_rx;
	schedule osdram_ba1 SB iuart0_rx;
	schedule osdram_cs SB iuart0_rx;
	schedule osdram_ras SB iuart0_rx;
	schedule osdram_cas SB iuart0_rx;
	schedule osdram_we SB iuart0_rx;
	schedule osdram_clk SB iuart0_rx;
	schedule osdram_cke SB iuart0_rx;
	schedule ospi1_ncs SB iuart0_rx;
	schedule ospi1_clk SB iuart0_rx;
	schedule ospi1_mosi SB iuart0_rx;
	schedule itms C itms;
	schedule itms CF itrst;
	schedule itms CF itck;
	schedule itms CF itdi;
	schedule itms CF ispi1_miso;
	schedule itms CF iboot_mode0;
	schedule itms CF iboot_mode1;
	schedule itms CF itest_mode;
	schedule ospi0_ncs SB itms;
	schedule ospi0_clk SB itms;
	schedule ospi0_mosi SB itms;
	schedule oqspi0_clk SB itms;
	schedule oqspi0_ncs SB itms;
	schedule ouart0_tx SB itms;
	schedule otdo SB itms;
	schedule osdram_a0 SB itms;
	schedule osdram_a1 SB itms;
	schedule osdram_a2 SB itms;
	schedule osdram_a3 SB itms;
	schedule osdram_a4 SB itms;
	schedule osdram_a5 SB itms;
	schedule osdram_a6 SB itms;
	schedule osdram_a7 SB itms;
	schedule osdram_a8 SB itms;
	schedule osdram_a9 SB itms;
	schedule osdram_a10 SB itms;
	schedule osdram_a11 SB itms;
	schedule osdram_a12 SB itms;
	schedule osdram_dq0 SB itms;
	schedule osdram_dq1 SB itms;
	schedule osdram_dq2 SB itms;
	schedule osdram_dq3 SB itms;
	schedule osdram_ba0 SB itms;
	schedule osdram_ba1 SB itms;
	schedule osdram_cs SB itms;
	schedule osdram_ras SB itms;
	schedule osdram_cas SB itms;
	schedule osdram_we SB itms;
	schedule osdram_clk SB itms;
	schedule osdram_cke SB itms;
	schedule ospi1_ncs SB itms;
	schedule ospi1_clk SB itms;
	schedule ospi1_mosi SB itms;
	schedule itrst C itrst;
	schedule itrst CF itck;
	schedule itrst CF itdi;
	schedule itrst CF ispi1_miso;
	schedule itrst CF iboot_mode0;
	schedule itrst CF iboot_mode1;
	schedule itrst CF itest_mode;
	schedule ospi0_ncs SB itrst;
	schedule ospi0_clk SB itrst;
	schedule ospi0_mosi SB itrst;
	schedule oqspi0_clk SB itrst;
	schedule oqspi0_ncs SB itrst;
	schedule ouart0_tx SB itrst;
	schedule otdo SB itrst;
	schedule osdram_a0 SB itrst;
	schedule osdram_a1 SB itrst;
	schedule osdram_a2 SB itrst;
	schedule osdram_a3 SB itrst;
	schedule osdram_a4 SB itrst;
	schedule osdram_a5 SB itrst;
	schedule osdram_a6 SB itrst;
	schedule osdram_a7 SB itrst;
	schedule osdram_a8 SB itrst;
	schedule osdram_a9 SB itrst;
	schedule osdram_a10 SB itrst;
	schedule osdram_a11 SB itrst;
	schedule osdram_a12 SB itrst;
	schedule osdram_dq0 SB itrst;
	schedule osdram_dq1 SB itrst;
	schedule osdram_dq2 SB itrst;
	schedule osdram_dq3 SB itrst;
	schedule osdram_ba0 SB itrst;
	schedule osdram_ba1 SB itrst;
	schedule osdram_cs SB itrst;
	schedule osdram_ras SB itrst;
	schedule osdram_cas SB itrst;
	schedule osdram_we SB itrst;
	schedule osdram_clk SB itrst;
	schedule osdram_cke SB itrst;
	schedule ospi1_ncs SB itrst;
	schedule ospi1_clk SB itrst;
	schedule ospi1_mosi SB itrst;
	schedule itck C itck;
	schedule itck CF itdi;
	schedule itck CF ispi1_miso;
	schedule itck CF iboot_mode0;
	schedule itck CF iboot_mode1;
	schedule itck CF itest_mode;
	schedule ospi0_ncs SB itck;
	schedule ospi0_clk SB itck;
	schedule ospi0_mosi SB itck;
	schedule oqspi0_clk SB itck;
	schedule oqspi0_ncs SB itck;
	schedule ouart0_tx SB itck;
	schedule otdo SB itck;
	schedule osdram_a0 SB itck;
	schedule osdram_a1 SB itck;
	schedule osdram_a2 SB itck;
	schedule osdram_a3 SB itck;
	schedule osdram_a4 SB itck;
	schedule osdram_a5 SB itck;
	schedule osdram_a6 SB itck;
	schedule osdram_a7 SB itck;
	schedule osdram_a8 SB itck;
	schedule osdram_a9 SB itck;
	schedule osdram_a10 SB itck;
	schedule osdram_a11 SB itck;
	schedule osdram_a12 SB itck;
	schedule osdram_dq0 SB itck;
	schedule osdram_dq1 SB itck;
	schedule osdram_dq2 SB itck;
	schedule osdram_dq3 SB itck;
	schedule osdram_ba0 SB itck;
	schedule osdram_ba1 SB itck;
	schedule osdram_cs SB itck;
	schedule osdram_ras SB itck;
	schedule osdram_cas SB itck;
	schedule osdram_we SB itck;
	schedule osdram_clk SB itck;
	schedule osdram_cke SB itck;
	schedule ospi1_ncs SB itck;
	schedule ospi1_clk SB itck;
	schedule ospi1_mosi SB itck;
	schedule itdi C itdi;
	schedule itdi CF ispi1_miso;
	schedule itdi CF iboot_mode0;
	schedule itdi CF iboot_mode1;
	schedule itdi CF itest_mode;
	schedule ospi0_ncs SB itdi;
	schedule ospi0_clk SB itdi;
	schedule ospi0_mosi SB itdi;
	schedule oqspi0_clk SB itdi;
	schedule oqspi0_ncs SB itdi;
	schedule ouart0_tx SB itdi;
	schedule otdo SB itdi;
	schedule osdram_a0 SB itdi;
	schedule osdram_a1 SB itdi;
	schedule osdram_a2 SB itdi;
	schedule osdram_a3 SB itdi;
	schedule osdram_a4 SB itdi;
	schedule osdram_a5 SB itdi;
	schedule osdram_a6 SB itdi;
	schedule osdram_a7 SB itdi;
	schedule osdram_a8 SB itdi;
	schedule osdram_a9 SB itdi;
	schedule osdram_a10 SB itdi;
	schedule osdram_a11 SB itdi;
	schedule osdram_a12 SB itdi;
	schedule osdram_dq0 SB itdi;
	schedule osdram_dq1 SB itdi;
	schedule osdram_dq2 SB itdi;
	schedule osdram_dq3 SB itdi;
	schedule osdram_ba0 SB itdi;
	schedule osdram_ba1 SB itdi;
	schedule osdram_cs SB itdi;
	schedule osdram_ras SB itdi;
	schedule osdram_cas SB itdi;
	schedule osdram_we SB itdi;
	schedule osdram_clk SB itdi;
	schedule osdram_cke SB itdi;
	schedule ospi1_ncs SB itdi;
	schedule ospi1_clk SB itdi;
	schedule ospi1_mosi SB itdi;
	schedule ispi1_miso C ispi1_miso;
	schedule ispi1_miso CF iboot_mode0;
	schedule ispi1_miso CF iboot_mode1;
	schedule ispi1_miso CF itest_mode;
	schedule ospi0_ncs SB ispi1_miso;
	schedule ospi0_clk SB ispi1_miso;
	schedule ospi0_mosi SB ispi1_miso;
	schedule oqspi0_clk SB ispi1_miso;
	schedule oqspi0_ncs SB ispi1_miso;
	schedule ouart0_tx SB ispi1_miso;
	schedule otdo SB ispi1_miso;
	schedule osdram_a0 SB ispi1_miso;
	schedule osdram_a1 SB ispi1_miso;
	schedule osdram_a2 SB ispi1_miso;
	schedule osdram_a3 SB ispi1_miso;
	schedule osdram_a4 SB ispi1_miso;
	schedule osdram_a5 SB ispi1_miso;
	schedule osdram_a6 SB ispi1_miso;
	schedule osdram_a7 SB ispi1_miso;
	schedule osdram_a8 SB ispi1_miso;
	schedule osdram_a9 SB ispi1_miso;
	schedule osdram_a10 SB ispi1_miso;
	schedule osdram_a11 SB ispi1_miso;
	schedule osdram_a12 SB ispi1_miso;
	schedule osdram_dq0 SB ispi1_miso;
	schedule osdram_dq1 SB ispi1_miso;
	schedule osdram_dq2 SB ispi1_miso;
	schedule osdram_dq3 SB ispi1_miso;
	schedule osdram_ba0 SB ispi1_miso;
	schedule osdram_ba1 SB ispi1_miso;
	schedule osdram_cs SB ispi1_miso;
	schedule osdram_ras SB ispi1_miso;
	schedule osdram_cas SB ispi1_miso;
	schedule osdram_we SB ispi1_miso;
	schedule osdram_clk SB ispi1_miso;
	schedule osdram_cke SB ispi1_miso;
	schedule ospi1_ncs SB ispi1_miso;
	schedule ospi1_clk SB ispi1_miso;
	schedule ospi1_mosi SB ispi1_miso;
	schedule iboot_mode0 C iboot_mode0;
	schedule iboot_mode0 CF iboot_mode1;
	schedule iboot_mode0 CF itest_mode;
	schedule ospi0_ncs SB iboot_mode0;
	schedule ospi0_clk SB iboot_mode0;
	schedule ospi0_mosi SB iboot_mode0;
	schedule oqspi0_clk SB iboot_mode0;
	schedule oqspi0_ncs SB iboot_mode0;
	schedule ouart0_tx SB iboot_mode0;
	schedule otdo SB iboot_mode0;
	schedule osdram_a0 SB iboot_mode0;
	schedule osdram_a1 SB iboot_mode0;
	schedule osdram_a2 SB iboot_mode0;
	schedule osdram_a3 SB iboot_mode0;
	schedule osdram_a4 SB iboot_mode0;
	schedule osdram_a5 SB iboot_mode0;
	schedule osdram_a6 SB iboot_mode0;
	schedule osdram_a7 SB iboot_mode0;
	schedule osdram_a8 SB iboot_mode0;
	schedule osdram_a9 SB iboot_mode0;
	schedule osdram_a10 SB iboot_mode0;
	schedule osdram_a11 SB iboot_mode0;
	schedule osdram_a12 SB iboot_mode0;
	schedule osdram_dq0 SB iboot_mode0;
	schedule osdram_dq1 SB iboot_mode0;
	schedule osdram_dq2 SB iboot_mode0;
	schedule osdram_dq3 SB iboot_mode0;
	schedule osdram_ba0 SB iboot_mode0;
	schedule osdram_ba1 SB iboot_mode0;
	schedule osdram_cs SB iboot_mode0;
	schedule osdram_ras SB iboot_mode0;
	schedule osdram_cas SB iboot_mode0;
	schedule osdram_we SB iboot_mode0;
	schedule osdram_clk SB iboot_mode0;
	schedule osdram_cke SB iboot_mode0;
	schedule ospi1_ncs SB iboot_mode0;
	schedule ospi1_clk SB iboot_mode0;
	schedule ospi1_mosi SB iboot_mode0;
	schedule iboot_mode1 C iboot_mode1;
	schedule iboot_mode1 CF itest_mode;
	schedule ospi0_ncs SB iboot_mode1;
	schedule ospi0_clk SB iboot_mode1;
	schedule ospi0_mosi SB iboot_mode1;
	schedule oqspi0_clk SB iboot_mode1;
	schedule oqspi0_ncs SB iboot_mode1;
	schedule ouart0_tx SB iboot_mode1;
	schedule otdo SB iboot_mode1;
	schedule osdram_a0 SB iboot_mode1;
	schedule osdram_a1 SB iboot_mode1;
	schedule osdram_a2 SB iboot_mode1;
	schedule osdram_a3 SB iboot_mode1;
	schedule osdram_a4 SB iboot_mode1;
	schedule osdram_a5 SB iboot_mode1;
	schedule osdram_a6 SB iboot_mode1;
	schedule osdram_a7 SB iboot_mode1;
	schedule osdram_a8 SB iboot_mode1;
	schedule osdram_a9 SB iboot_mode1;
	schedule osdram_a10 SB iboot_mode1;
	schedule osdram_a11 SB iboot_mode1;
	schedule osdram_a12 SB iboot_mode1;
	schedule osdram_dq0 SB iboot_mode1;
	schedule osdram_dq1 SB iboot_mode1;
	schedule osdram_dq2 SB iboot_mode1;
	schedule osdram_dq3 SB iboot_mode1;
	schedule osdram_ba0 SB iboot_mode1;
	schedule osdram_ba1 SB iboot_mode1;
	schedule osdram_cs SB iboot_mode1;
	schedule osdram_ras SB iboot_mode1;
	schedule osdram_cas SB iboot_mode1;
	schedule osdram_we SB iboot_mode1;
	schedule osdram_clk SB iboot_mode1;
	schedule osdram_cke SB iboot_mode1;
	schedule ospi1_ncs SB iboot_mode1;
	schedule ospi1_clk SB iboot_mode1;
	schedule ospi1_mosi SB iboot_mode1;
	schedule itest_mode C itest_mode;
	schedule ospi0_ncs SB itest_mode;
	schedule ospi0_clk SB itest_mode;
	schedule ospi0_mosi SB itest_mode;
	schedule oqspi0_clk SB itest_mode;
	schedule oqspi0_ncs SB itest_mode;
	schedule ouart0_tx SB itest_mode;
	schedule otdo SB itest_mode;
	schedule osdram_a0 SB itest_mode;
	schedule osdram_a1 SB itest_mode;
	schedule osdram_a2 SB itest_mode;
	schedule osdram_a3 SB itest_mode;
	schedule osdram_a4 SB itest_mode;
	schedule osdram_a5 SB itest_mode;
	schedule osdram_a6 SB itest_mode;
	schedule osdram_a7 SB itest_mode;
	schedule osdram_a8 SB itest_mode;
	schedule osdram_a9 SB itest_mode;
	schedule osdram_a10 SB itest_mode;
	schedule osdram_a11 SB itest_mode;
	schedule osdram_a12 SB itest_mode;
	schedule osdram_dq0 SB itest_mode;
	schedule osdram_dq1 SB itest_mode;
	schedule osdram_dq2 SB itest_mode;
	schedule osdram_dq3 SB itest_mode;
	schedule osdram_ba0 SB itest_mode;
	schedule osdram_ba1 SB itest_mode;
	schedule osdram_cs SB itest_mode;
	schedule osdram_ras SB itest_mode;
	schedule osdram_cas SB itest_mode;
	schedule osdram_we SB itest_mode;
	schedule osdram_clk SB itest_mode;
	schedule osdram_cke SB itest_mode;
	schedule ospi1_ncs SB itest_mode;
	schedule ospi1_clk SB itest_mode;
	schedule ospi1_mosi SB itest_mode;
	schedule ospi0_ncs CF ospi0_ncs;
	schedule ospi0_ncs CF ospi0_clk;
	schedule ospi0_ncs CF ospi0_mosi;
	schedule ospi0_ncs CF oqspi0_clk;
	schedule ospi0_ncs CF oqspi0_ncs;
	schedule ospi0_ncs CF ouart0_tx;
	schedule ospi0_ncs CF otdo;
	schedule ospi0_ncs CF osdram_a0;
	schedule ospi0_ncs CF osdram_a1;
	schedule ospi0_ncs CF osdram_a2;
	schedule ospi0_ncs CF osdram_a3;
	schedule ospi0_ncs CF osdram_a4;
	schedule ospi0_ncs CF osdram_a5;
	schedule ospi0_ncs CF osdram_a6;
	schedule ospi0_ncs CF osdram_a7;
	schedule ospi0_ncs CF osdram_a8;
	schedule ospi0_ncs CF osdram_a9;
	schedule ospi0_ncs CF osdram_a10;
	schedule ospi0_ncs CF osdram_a11;
	schedule ospi0_ncs CF osdram_a12;
	schedule ospi0_ncs CF osdram_dq0;
	schedule ospi0_ncs CF osdram_dq1;
	schedule ospi0_ncs CF osdram_dq2;
	schedule ospi0_ncs CF osdram_dq3;
	schedule ospi0_ncs CF osdram_ba0;
	schedule ospi0_ncs CF osdram_ba1;
	schedule ospi0_ncs CF osdram_cs;
	schedule ospi0_ncs CF osdram_ras;
	schedule ospi0_ncs CF osdram_cas;
	schedule ospi0_ncs CF osdram_we;
	schedule ospi0_ncs CF osdram_clk;
	schedule ospi0_ncs CF osdram_cke;
	schedule ospi0_ncs CF ospi1_ncs;
	schedule ospi0_ncs CF ospi1_clk;
	schedule ospi0_ncs CF ospi1_mosi;
	schedule ospi0_clk CF ospi0_clk;
	schedule ospi0_clk CF ospi0_mosi;
	schedule ospi0_clk CF oqspi0_clk;
	schedule ospi0_clk CF oqspi0_ncs;
	schedule ospi0_clk CF ouart0_tx;
	schedule ospi0_clk CF otdo;
	schedule ospi0_clk CF osdram_a0;
	schedule ospi0_clk CF osdram_a1;
	schedule ospi0_clk CF osdram_a2;
	schedule ospi0_clk CF osdram_a3;
	schedule ospi0_clk CF osdram_a4;
	schedule ospi0_clk CF osdram_a5;
	schedule ospi0_clk CF osdram_a6;
	schedule ospi0_clk CF osdram_a7;
	schedule ospi0_clk CF osdram_a8;
	schedule ospi0_clk CF osdram_a9;
	schedule ospi0_clk CF osdram_a10;
	schedule ospi0_clk CF osdram_a11;
	schedule ospi0_clk CF osdram_a12;
	schedule ospi0_clk CF osdram_dq0;
	schedule ospi0_clk CF osdram_dq1;
	schedule ospi0_clk CF osdram_dq2;
	schedule ospi0_clk CF osdram_dq3;
	schedule ospi0_clk CF osdram_ba0;
	schedule ospi0_clk CF osdram_ba1;
	schedule ospi0_clk CF osdram_cs;
	schedule ospi0_clk CF osdram_ras;
	schedule ospi0_clk CF osdram_cas;
	schedule ospi0_clk CF osdram_we;
	schedule ospi0_clk CF osdram_clk;
	schedule ospi0_clk CF osdram_cke;
	schedule ospi0_clk CF ospi1_ncs;
	schedule ospi0_clk CF ospi1_clk;
	schedule ospi0_clk CF ospi1_mosi;
	schedule ospi0_mosi CF ospi0_mosi;
	schedule ospi0_mosi CF oqspi0_clk;
	schedule ospi0_mosi CF oqspi0_ncs;
	schedule ospi0_mosi CF ouart0_tx;
	schedule ospi0_mosi CF otdo;
	schedule ospi0_mosi CF osdram_a0;
	schedule ospi0_mosi CF osdram_a1;
	schedule ospi0_mosi CF osdram_a2;
	schedule ospi0_mosi CF osdram_a3;
	schedule ospi0_mosi CF osdram_a4;
	schedule ospi0_mosi CF osdram_a5;
	schedule ospi0_mosi CF osdram_a6;
	schedule ospi0_mosi CF osdram_a7;
	schedule ospi0_mosi CF osdram_a8;
	schedule ospi0_mosi CF osdram_a9;
	schedule ospi0_mosi CF osdram_a10;
	schedule ospi0_mosi CF osdram_a11;
	schedule ospi0_mosi CF osdram_a12;
	schedule ospi0_mosi CF osdram_dq0;
	schedule ospi0_mosi CF osdram_dq1;
	schedule ospi0_mosi CF osdram_dq2;
	schedule ospi0_mosi CF osdram_dq3;
	schedule ospi0_mosi CF osdram_ba0;
	schedule ospi0_mosi CF osdram_ba1;
	schedule ospi0_mosi CF osdram_cs;
	schedule ospi0_mosi CF osdram_ras;
	schedule ospi0_mosi CF osdram_cas;
	schedule ospi0_mosi CF osdram_we;
	schedule ospi0_mosi CF osdram_clk;
	schedule ospi0_mosi CF osdram_cke;
	schedule ospi0_mosi CF ospi1_ncs;
	schedule ospi0_mosi CF ospi1_clk;
	schedule ospi0_mosi CF ospi1_mosi;
	schedule oqspi0_clk CF oqspi0_clk;
	schedule oqspi0_clk CF oqspi0_ncs;
	schedule oqspi0_clk CF ouart0_tx;
	schedule oqspi0_clk CF otdo;
	schedule oqspi0_clk CF osdram_a0;
	schedule oqspi0_clk CF osdram_a1;
	schedule oqspi0_clk CF osdram_a2;
	schedule oqspi0_clk CF osdram_a3;
	schedule oqspi0_clk CF osdram_a4;
	schedule oqspi0_clk CF osdram_a5;
	schedule oqspi0_clk CF osdram_a6;
	schedule oqspi0_clk CF osdram_a7;
	schedule oqspi0_clk CF osdram_a8;
	schedule oqspi0_clk CF osdram_a9;
	schedule oqspi0_clk CF osdram_a10;
	schedule oqspi0_clk CF osdram_a11;
	schedule oqspi0_clk CF osdram_a12;
	schedule oqspi0_clk CF osdram_dq0;
	schedule oqspi0_clk CF osdram_dq1;
	schedule oqspi0_clk CF osdram_dq2;
	schedule oqspi0_clk CF osdram_dq3;
	schedule oqspi0_clk CF osdram_ba0;
	schedule oqspi0_clk CF osdram_ba1;
	schedule oqspi0_clk CF osdram_cs;
	schedule oqspi0_clk CF osdram_ras;
	schedule oqspi0_clk CF osdram_cas;
	schedule oqspi0_clk CF osdram_we;
	schedule oqspi0_clk CF osdram_clk;
	schedule oqspi0_clk CF osdram_cke;
	schedule oqspi0_clk CF ospi1_ncs;
	schedule oqspi0_clk CF ospi1_clk;
	schedule oqspi0_clk CF ospi1_mosi;
	schedule oqspi0_ncs CF oqspi0_ncs;
	schedule oqspi0_ncs CF ouart0_tx;
	schedule oqspi0_ncs CF otdo;
	schedule oqspi0_ncs CF osdram_a0;
	schedule oqspi0_ncs CF osdram_a1;
	schedule oqspi0_ncs CF osdram_a2;
	schedule oqspi0_ncs CF osdram_a3;
	schedule oqspi0_ncs CF osdram_a4;
	schedule oqspi0_ncs CF osdram_a5;
	schedule oqspi0_ncs CF osdram_a6;
	schedule oqspi0_ncs CF osdram_a7;
	schedule oqspi0_ncs CF osdram_a8;
	schedule oqspi0_ncs CF osdram_a9;
	schedule oqspi0_ncs CF osdram_a10;
	schedule oqspi0_ncs CF osdram_a11;
	schedule oqspi0_ncs CF osdram_a12;
	schedule oqspi0_ncs CF osdram_dq0;
	schedule oqspi0_ncs CF osdram_dq1;
	schedule oqspi0_ncs CF osdram_dq2;
	schedule oqspi0_ncs CF osdram_dq3;
	schedule oqspi0_ncs CF osdram_ba0;
	schedule oqspi0_ncs CF osdram_ba1;
	schedule oqspi0_ncs CF osdram_cs;
	schedule oqspi0_ncs CF osdram_ras;
	schedule oqspi0_ncs CF osdram_cas;
	schedule oqspi0_ncs CF osdram_we;
	schedule oqspi0_ncs CF osdram_clk;
	schedule oqspi0_ncs CF osdram_cke;
	schedule oqspi0_ncs CF ospi1_ncs;
	schedule oqspi0_ncs CF ospi1_clk;
	schedule oqspi0_ncs CF ospi1_mosi;
	schedule ouart0_tx CF ouart0_tx;
	schedule ouart0_tx CF otdo;
	schedule ouart0_tx CF osdram_a0;
	schedule ouart0_tx CF osdram_a1;
	schedule ouart0_tx CF osdram_a2;
	schedule ouart0_tx CF osdram_a3;
	schedule ouart0_tx CF osdram_a4;
	schedule ouart0_tx CF osdram_a5;
	schedule ouart0_tx CF osdram_a6;
	schedule ouart0_tx CF osdram_a7;
	schedule ouart0_tx CF osdram_a8;
	schedule ouart0_tx CF osdram_a9;
	schedule ouart0_tx CF osdram_a10;
	schedule ouart0_tx CF osdram_a11;
	schedule ouart0_tx CF osdram_a12;
	schedule ouart0_tx CF osdram_dq0;
	schedule ouart0_tx CF osdram_dq1;
	schedule ouart0_tx CF osdram_dq2;
	schedule ouart0_tx CF osdram_dq3;
	schedule ouart0_tx CF osdram_ba0;
	schedule ouart0_tx CF osdram_ba1;
	schedule ouart0_tx CF osdram_cs;
	schedule ouart0_tx CF osdram_ras;
	schedule ouart0_tx CF osdram_cas;
	schedule ouart0_tx CF osdram_we;
	schedule ouart0_tx CF osdram_clk;
	schedule ouart0_tx CF osdram_cke;
	schedule ouart0_tx CF ospi1_ncs;
	schedule ouart0_tx CF ospi1_clk;
	schedule ouart0_tx CF ospi1_mosi;
	schedule otdo CF otdo;
	schedule otdo CF osdram_a0;
	schedule otdo CF osdram_a1;
	schedule otdo CF osdram_a2;
	schedule otdo CF osdram_a3;
	schedule otdo CF osdram_a4;
	schedule otdo CF osdram_a5;
	schedule otdo CF osdram_a6;
	schedule otdo CF osdram_a7;
	schedule otdo CF osdram_a8;
	schedule otdo CF osdram_a9;
	schedule otdo CF osdram_a10;
	schedule otdo CF osdram_a11;
	schedule otdo CF osdram_a12;
	schedule otdo CF osdram_dq0;
	schedule otdo CF osdram_dq1;
	schedule otdo CF osdram_dq2;
	schedule otdo CF osdram_dq3;
	schedule otdo CF osdram_ba0;
	schedule otdo CF osdram_ba1;
	schedule otdo CF osdram_cs;
	schedule otdo CF osdram_ras;
	schedule otdo CF osdram_cas;
	schedule otdo CF osdram_we;
	schedule otdo CF osdram_clk;
	schedule otdo CF osdram_cke;
	schedule otdo CF ospi1_ncs;
	schedule otdo CF ospi1_clk;
	schedule otdo CF ospi1_mosi;
	schedule osdram_a0 CF osdram_a0;
	schedule osdram_a0 CF osdram_a1;
	schedule osdram_a0 CF osdram_a2;
	schedule osdram_a0 CF osdram_a3;
	schedule osdram_a0 CF osdram_a4;
	schedule osdram_a0 CF osdram_a5;
	schedule osdram_a0 CF osdram_a6;
	schedule osdram_a0 CF osdram_a7;
	schedule osdram_a0 CF osdram_a8;
	schedule osdram_a0 CF osdram_a9;
	schedule osdram_a0 CF osdram_a10;
	schedule osdram_a0 CF osdram_a11;
	schedule osdram_a0 CF osdram_a12;
	schedule osdram_a0 CF osdram_dq0;
	schedule osdram_a0 CF osdram_dq1;
	schedule osdram_a0 CF osdram_dq2;
	schedule osdram_a0 CF osdram_dq3;
	schedule osdram_a0 CF osdram_ba0;
	schedule osdram_a0 CF osdram_ba1;
	schedule osdram_a0 CF osdram_cs;
	schedule osdram_a0 CF osdram_ras;
	schedule osdram_a0 CF osdram_cas;
	schedule osdram_a0 CF osdram_we;
	schedule osdram_a0 CF osdram_clk;
	schedule osdram_a0 CF osdram_cke;
	schedule osdram_a0 CF ospi1_ncs;
	schedule osdram_a0 CF ospi1_clk;
	schedule osdram_a0 CF ospi1_mosi;
	schedule osdram_a1 CF osdram_a1;
	schedule osdram_a1 CF osdram_a2;
	schedule osdram_a1 CF osdram_a3;
	schedule osdram_a1 CF osdram_a4;
	schedule osdram_a1 CF osdram_a5;
	schedule osdram_a1 CF osdram_a6;
	schedule osdram_a1 CF osdram_a7;
	schedule osdram_a1 CF osdram_a8;
	schedule osdram_a1 CF osdram_a9;
	schedule osdram_a1 CF osdram_a10;
	schedule osdram_a1 CF osdram_a11;
	schedule osdram_a1 CF osdram_a12;
	schedule osdram_a1 CF osdram_dq0;
	schedule osdram_a1 CF osdram_dq1;
	schedule osdram_a1 CF osdram_dq2;
	schedule osdram_a1 CF osdram_dq3;
	schedule osdram_a1 CF osdram_ba0;
	schedule osdram_a1 CF osdram_ba1;
	schedule osdram_a1 CF osdram_cs;
	schedule osdram_a1 CF osdram_ras;
	schedule osdram_a1 CF osdram_cas;
	schedule osdram_a1 CF osdram_we;
	schedule osdram_a1 CF osdram_clk;
	schedule osdram_a1 CF osdram_cke;
	schedule osdram_a1 CF ospi1_ncs;
	schedule osdram_a1 CF ospi1_clk;
	schedule osdram_a1 CF ospi1_mosi;
	schedule osdram_a2 CF osdram_a2;
	schedule osdram_a2 CF osdram_a3;
	schedule osdram_a2 CF osdram_a4;
	schedule osdram_a2 CF osdram_a5;
	schedule osdram_a2 CF osdram_a6;
	schedule osdram_a2 CF osdram_a7;
	schedule osdram_a2 CF osdram_a8;
	schedule osdram_a2 CF osdram_a9;
	schedule osdram_a2 CF osdram_a10;
	schedule osdram_a2 CF osdram_a11;
	schedule osdram_a2 CF osdram_a12;
	schedule osdram_a2 CF osdram_dq0;
	schedule osdram_a2 CF osdram_dq1;
	schedule osdram_a2 CF osdram_dq2;
	schedule osdram_a2 CF osdram_dq3;
	schedule osdram_a2 CF osdram_ba0;
	schedule osdram_a2 CF osdram_ba1;
	schedule osdram_a2 CF osdram_cs;
	schedule osdram_a2 CF osdram_ras;
	schedule osdram_a2 CF osdram_cas;
	schedule osdram_a2 CF osdram_we;
	schedule osdram_a2 CF osdram_clk;
	schedule osdram_a2 CF osdram_cke;
	schedule osdram_a2 CF ospi1_ncs;
	schedule osdram_a2 CF ospi1_clk;
	schedule osdram_a2 CF ospi1_mosi;
	schedule osdram_a3 CF osdram_a3;
	schedule osdram_a3 CF osdram_a4;
	schedule osdram_a3 CF osdram_a5;
	schedule osdram_a3 CF osdram_a6;
	schedule osdram_a3 CF osdram_a7;
	schedule osdram_a3 CF osdram_a8;
	schedule osdram_a3 CF osdram_a9;
	schedule osdram_a3 CF osdram_a10;
	schedule osdram_a3 CF osdram_a11;
	schedule osdram_a3 CF osdram_a12;
	schedule osdram_a3 CF osdram_dq0;
	schedule osdram_a3 CF osdram_dq1;
	schedule osdram_a3 CF osdram_dq2;
	schedule osdram_a3 CF osdram_dq3;
	schedule osdram_a3 CF osdram_ba0;
	schedule osdram_a3 CF osdram_ba1;
	schedule osdram_a3 CF osdram_cs;
	schedule osdram_a3 CF osdram_ras;
	schedule osdram_a3 CF osdram_cas;
	schedule osdram_a3 CF osdram_we;
	schedule osdram_a3 CF osdram_clk;
	schedule osdram_a3 CF osdram_cke;
	schedule osdram_a3 CF ospi1_ncs;
	schedule osdram_a3 CF ospi1_clk;
	schedule osdram_a3 CF ospi1_mosi;
	schedule osdram_a4 CF osdram_a4;
	schedule osdram_a4 CF osdram_a5;
	schedule osdram_a4 CF osdram_a6;
	schedule osdram_a4 CF osdram_a7;
	schedule osdram_a4 CF osdram_a8;
	schedule osdram_a4 CF osdram_a9;
	schedule osdram_a4 CF osdram_a10;
	schedule osdram_a4 CF osdram_a11;
	schedule osdram_a4 CF osdram_a12;
	schedule osdram_a4 CF osdram_dq0;
	schedule osdram_a4 CF osdram_dq1;
	schedule osdram_a4 CF osdram_dq2;
	schedule osdram_a4 CF osdram_dq3;
	schedule osdram_a4 CF osdram_ba0;
	schedule osdram_a4 CF osdram_ba1;
	schedule osdram_a4 CF osdram_cs;
	schedule osdram_a4 CF osdram_ras;
	schedule osdram_a4 CF osdram_cas;
	schedule osdram_a4 CF osdram_we;
	schedule osdram_a4 CF osdram_clk;
	schedule osdram_a4 CF osdram_cke;
	schedule osdram_a4 CF ospi1_ncs;
	schedule osdram_a4 CF ospi1_clk;
	schedule osdram_a4 CF ospi1_mosi;
	schedule osdram_a5 CF osdram_a5;
	schedule osdram_a5 CF osdram_a6;
	schedule osdram_a5 CF osdram_a7;
	schedule osdram_a5 CF osdram_a8;
	schedule osdram_a5 CF osdram_a9;
	schedule osdram_a5 CF osdram_a10;
	schedule osdram_a5 CF osdram_a11;
	schedule osdram_a5 CF osdram_a12;
	schedule osdram_a5 CF osdram_dq0;
	schedule osdram_a5 CF osdram_dq1;
	schedule osdram_a5 CF osdram_dq2;
	schedule osdram_a5 CF osdram_dq3;
	schedule osdram_a5 CF osdram_ba0;
	schedule osdram_a5 CF osdram_ba1;
	schedule osdram_a5 CF osdram_cs;
	schedule osdram_a5 CF osdram_ras;
	schedule osdram_a5 CF osdram_cas;
	schedule osdram_a5 CF osdram_we;
	schedule osdram_a5 CF osdram_clk;
	schedule osdram_a5 CF osdram_cke;
	schedule osdram_a5 CF ospi1_ncs;
	schedule osdram_a5 CF ospi1_clk;
	schedule osdram_a5 CF ospi1_mosi;
	schedule osdram_a6 CF osdram_a6;
	schedule osdram_a6 CF osdram_a7;
	schedule osdram_a6 CF osdram_a8;
	schedule osdram_a6 CF osdram_a9;
	schedule osdram_a6 CF osdram_a10;
	schedule osdram_a6 CF osdram_a11;
	schedule osdram_a6 CF osdram_a12;
	schedule osdram_a6 CF osdram_dq0;
	schedule osdram_a6 CF osdram_dq1;
	schedule osdram_a6 CF osdram_dq2;
	schedule osdram_a6 CF osdram_dq3;
	schedule osdram_a6 CF osdram_ba0;
	schedule osdram_a6 CF osdram_ba1;
	schedule osdram_a6 CF osdram_cs;
	schedule osdram_a6 CF osdram_ras;
	schedule osdram_a6 CF osdram_cas;
	schedule osdram_a6 CF osdram_we;
	schedule osdram_a6 CF osdram_clk;
	schedule osdram_a6 CF osdram_cke;
	schedule osdram_a6 CF ospi1_ncs;
	schedule osdram_a6 CF ospi1_clk;
	schedule osdram_a6 CF ospi1_mosi;
	schedule osdram_a7 CF osdram_a7;
	schedule osdram_a7 CF osdram_a8;
	schedule osdram_a7 CF osdram_a9;
	schedule osdram_a7 CF osdram_a10;
	schedule osdram_a7 CF osdram_a11;
	schedule osdram_a7 CF osdram_a12;
	schedule osdram_a7 CF osdram_dq0;
	schedule osdram_a7 CF osdram_dq1;
	schedule osdram_a7 CF osdram_dq2;
	schedule osdram_a7 CF osdram_dq3;
	schedule osdram_a7 CF osdram_ba0;
	schedule osdram_a7 CF osdram_ba1;
	schedule osdram_a7 CF osdram_cs;
	schedule osdram_a7 CF osdram_ras;
	schedule osdram_a7 CF osdram_cas;
	schedule osdram_a7 CF osdram_we;
	schedule osdram_a7 CF osdram_clk;
	schedule osdram_a7 CF osdram_cke;
	schedule osdram_a7 CF ospi1_ncs;
	schedule osdram_a7 CF ospi1_clk;
	schedule osdram_a7 CF ospi1_mosi;
	schedule osdram_a8 CF osdram_a8;
	schedule osdram_a8 CF osdram_a9;
	schedule osdram_a8 CF osdram_a10;
	schedule osdram_a8 CF osdram_a11;
	schedule osdram_a8 CF osdram_a12;
	schedule osdram_a8 CF osdram_dq0;
	schedule osdram_a8 CF osdram_dq1;
	schedule osdram_a8 CF osdram_dq2;
	schedule osdram_a8 CF osdram_dq3;
	schedule osdram_a8 CF osdram_ba0;
	schedule osdram_a8 CF osdram_ba1;
	schedule osdram_a8 CF osdram_cs;
	schedule osdram_a8 CF osdram_ras;
	schedule osdram_a8 CF osdram_cas;
	schedule osdram_a8 CF osdram_we;
	schedule osdram_a8 CF osdram_clk;
	schedule osdram_a8 CF osdram_cke;
	schedule osdram_a8 CF ospi1_ncs;
	schedule osdram_a8 CF ospi1_clk;
	schedule osdram_a8 CF ospi1_mosi;
	schedule osdram_a9 CF osdram_a9;
	schedule osdram_a9 CF osdram_a10;
	schedule osdram_a9 CF osdram_a11;
	schedule osdram_a9 CF osdram_a12;
	schedule osdram_a9 CF osdram_dq0;
	schedule osdram_a9 CF osdram_dq1;
	schedule osdram_a9 CF osdram_dq2;
	schedule osdram_a9 CF osdram_dq3;
	schedule osdram_a9 CF osdram_ba0;
	schedule osdram_a9 CF osdram_ba1;
	schedule osdram_a9 CF osdram_cs;
	schedule osdram_a9 CF osdram_ras;
	schedule osdram_a9 CF osdram_cas;
	schedule osdram_a9 CF osdram_we;
	schedule osdram_a9 CF osdram_clk;
	schedule osdram_a9 CF osdram_cke;
	schedule osdram_a9 CF ospi1_ncs;
	schedule osdram_a9 CF ospi1_clk;
	schedule osdram_a9 CF ospi1_mosi;
	schedule osdram_a10 CF osdram_a10;
	schedule osdram_a10 CF osdram_a11;
	schedule osdram_a10 CF osdram_a12;
	schedule osdram_a10 CF osdram_dq0;
	schedule osdram_a10 CF osdram_dq1;
	schedule osdram_a10 CF osdram_dq2;
	schedule osdram_a10 CF osdram_dq3;
	schedule osdram_a10 CF osdram_ba0;
	schedule osdram_a10 CF osdram_ba1;
	schedule osdram_a10 CF osdram_cs;
	schedule osdram_a10 CF osdram_ras;
	schedule osdram_a10 CF osdram_cas;
	schedule osdram_a10 CF osdram_we;
	schedule osdram_a10 CF osdram_clk;
	schedule osdram_a10 CF osdram_cke;
	schedule osdram_a10 CF ospi1_ncs;
	schedule osdram_a10 CF ospi1_clk;
	schedule osdram_a10 CF ospi1_mosi;
	schedule osdram_a11 CF osdram_a11;
	schedule osdram_a11 CF osdram_a12;
	schedule osdram_a11 CF osdram_dq0;
	schedule osdram_a11 CF osdram_dq1;
	schedule osdram_a11 CF osdram_dq2;
	schedule osdram_a11 CF osdram_dq3;
	schedule osdram_a11 CF osdram_ba0;
	schedule osdram_a11 CF osdram_ba1;
	schedule osdram_a11 CF osdram_cs;
	schedule osdram_a11 CF osdram_ras;
	schedule osdram_a11 CF osdram_cas;
	schedule osdram_a11 CF osdram_we;
	schedule osdram_a11 CF osdram_clk;
	schedule osdram_a11 CF osdram_cke;
	schedule osdram_a11 CF ospi1_ncs;
	schedule osdram_a11 CF ospi1_clk;
	schedule osdram_a11 CF ospi1_mosi;
	schedule osdram_a12 CF osdram_a12;
	schedule osdram_a12 CF osdram_dq0;
	schedule osdram_a12 CF osdram_dq1;
	schedule osdram_a12 CF osdram_dq2;
	schedule osdram_a12 CF osdram_dq3;
	schedule osdram_a12 CF osdram_ba0;
	schedule osdram_a12 CF osdram_ba1;
	schedule osdram_a12 CF osdram_cs;
	schedule osdram_a12 CF osdram_ras;
	schedule osdram_a12 CF osdram_cas;
	schedule osdram_a12 CF osdram_we;
	schedule osdram_a12 CF osdram_clk;
	schedule osdram_a12 CF osdram_cke;
	schedule osdram_a12 CF ospi1_ncs;
	schedule osdram_a12 CF ospi1_clk;
	schedule osdram_a12 CF ospi1_mosi;
	schedule osdram_dq0 CF osdram_dq0;
	schedule osdram_dq0 CF osdram_dq1;
	schedule osdram_dq0 CF osdram_dq2;
	schedule osdram_dq0 CF osdram_dq3;
	schedule osdram_dq0 CF osdram_ba0;
	schedule osdram_dq0 CF osdram_ba1;
	schedule osdram_dq0 CF osdram_cs;
	schedule osdram_dq0 CF osdram_ras;
	schedule osdram_dq0 CF osdram_cas;
	schedule osdram_dq0 CF osdram_we;
	schedule osdram_dq0 CF osdram_clk;
	schedule osdram_dq0 CF osdram_cke;
	schedule osdram_dq0 CF ospi1_ncs;
	schedule osdram_dq0 CF ospi1_clk;
	schedule osdram_dq0 CF ospi1_mosi;
	schedule osdram_dq1 CF osdram_dq1;
	schedule osdram_dq1 CF osdram_dq2;
	schedule osdram_dq1 CF osdram_dq3;
	schedule osdram_dq1 CF osdram_ba0;
	schedule osdram_dq1 CF osdram_ba1;
	schedule osdram_dq1 CF osdram_cs;
	schedule osdram_dq1 CF osdram_ras;
	schedule osdram_dq1 CF osdram_cas;
	schedule osdram_dq1 CF osdram_we;
	schedule osdram_dq1 CF osdram_clk;
	schedule osdram_dq1 CF osdram_cke;
	schedule osdram_dq1 CF ospi1_ncs;
	schedule osdram_dq1 CF ospi1_clk;
	schedule osdram_dq1 CF ospi1_mosi;
	schedule osdram_dq2 CF osdram_dq2;
	schedule osdram_dq2 CF osdram_dq3;
	schedule osdram_dq2 CF osdram_ba0;
	schedule osdram_dq2 CF osdram_ba1;
	schedule osdram_dq2 CF osdram_cs;
	schedule osdram_dq2 CF osdram_ras;
	schedule osdram_dq2 CF osdram_cas;
	schedule osdram_dq2 CF osdram_we;
	schedule osdram_dq2 CF osdram_clk;
	schedule osdram_dq2 CF osdram_cke;
	schedule osdram_dq2 CF ospi1_ncs;
	schedule osdram_dq2 CF ospi1_clk;
	schedule osdram_dq2 CF ospi1_mosi;
	schedule osdram_dq3 CF osdram_dq3;
	schedule osdram_dq3 CF osdram_ba0;
	schedule osdram_dq3 CF osdram_ba1;
	schedule osdram_dq3 CF osdram_cs;
	schedule osdram_dq3 CF osdram_ras;
	schedule osdram_dq3 CF osdram_cas;
	schedule osdram_dq3 CF osdram_we;
	schedule osdram_dq3 CF osdram_clk;
	schedule osdram_dq3 CF osdram_cke;
	schedule osdram_dq3 CF ospi1_ncs;
	schedule osdram_dq3 CF ospi1_clk;
	schedule osdram_dq3 CF ospi1_mosi;
	schedule osdram_ba0 CF osdram_ba0;
	schedule osdram_ba0 CF osdram_ba1;
	schedule osdram_ba0 CF osdram_cs;
	schedule osdram_ba0 CF osdram_ras;
	schedule osdram_ba0 CF osdram_cas;
	schedule osdram_ba0 CF osdram_we;
	schedule osdram_ba0 CF osdram_clk;
	schedule osdram_ba0 CF osdram_cke;
	schedule osdram_ba0 CF ospi1_ncs;
	schedule osdram_ba0 CF ospi1_clk;
	schedule osdram_ba0 CF ospi1_mosi;
	schedule osdram_ba1 CF osdram_ba1;
	schedule osdram_ba1 CF osdram_cs;
	schedule osdram_ba1 CF osdram_ras;
	schedule osdram_ba1 CF osdram_cas;
	schedule osdram_ba1 CF osdram_we;
	schedule osdram_ba1 CF osdram_clk;
	schedule osdram_ba1 CF osdram_cke;
	schedule osdram_ba1 CF ospi1_ncs;
	schedule osdram_ba1 CF ospi1_clk;
	schedule osdram_ba1 CF ospi1_mosi;
	schedule osdram_cs CF osdram_cs;
	schedule osdram_cs CF osdram_ras;
	schedule osdram_cs CF osdram_cas;
	schedule osdram_cs CF osdram_we;
	schedule osdram_cs CF osdram_clk;
	schedule osdram_cs CF osdram_cke;
	schedule osdram_cs CF ospi1_ncs;
	schedule osdram_cs CF ospi1_clk;
	schedule osdram_cs CF ospi1_mosi;
	schedule osdram_ras CF osdram_ras;
	schedule osdram_ras CF osdram_cas;
	schedule osdram_ras CF osdram_we;
	schedule osdram_ras CF osdram_clk;
	schedule osdram_ras CF osdram_cke;
	schedule osdram_ras CF ospi1_ncs;
	schedule osdram_ras CF ospi1_clk;
	schedule osdram_ras CF ospi1_mosi;
	schedule osdram_cas CF osdram_cas;
	schedule osdram_cas CF osdram_we;
	schedule osdram_cas CF osdram_clk;
	schedule osdram_cas CF osdram_cke;
	schedule osdram_cas CF ospi1_ncs;
	schedule osdram_cas CF ospi1_clk;
	schedule osdram_cas CF ospi1_mosi;
	schedule osdram_we CF osdram_we;
	schedule osdram_we CF osdram_clk;
	schedule osdram_we CF osdram_cke;
	schedule osdram_we CF ospi1_ncs;
	schedule osdram_we CF ospi1_clk;
	schedule osdram_we CF ospi1_mosi;
	schedule osdram_clk CF osdram_clk;
	schedule osdram_clk CF osdram_cke;
	schedule osdram_clk CF ospi1_ncs;
	schedule osdram_clk CF ospi1_clk;
	schedule osdram_clk CF ospi1_mosi;
	schedule osdram_cke CF osdram_cke;
	schedule osdram_cke CF ospi1_ncs;
	schedule osdram_cke CF ospi1_clk;
	schedule osdram_cke CF ospi1_mosi;
	schedule ospi1_ncs CF ospi1_ncs;
	schedule ospi1_ncs CF ospi1_clk;
	schedule ospi1_ncs CF ospi1_mosi;
	schedule ospi1_clk CF ospi1_clk;
	schedule ospi1_clk CF ospi1_mosi;
	schedule ospi1_mosi CF ospi1_mosi;
endmodule


