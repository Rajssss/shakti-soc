// Bluespec wrapper, created by Import BVI Wizard
// Created on: Wed Dec 04 13:11:05 IST 2019
// Created by: Sadhana
// Bluespec version: 2019.05.beta2 2019-05-24 a88bf40db


interface Ifc_aardonyx_wrapper;
	interface Inout#(Bit#(1)) ioGPIO_0;
	interface Inout#(Bit#(1)) ioGPIO_1;
	interface Inout#(Bit#(1)) ioGPIO_2;
	interface Inout#(Bit#(1)) ioGPIO_3;
	interface Inout#(Bit#(1)) ioGPIO_4;
	interface Inout#(Bit#(1)) ioGPIO_5;
	interface Inout#(Bit#(1)) ioGPIO_6;
	interface Inout#(Bit#(1)) ioGPIO_7;
	interface Inout#(Bit#(1)) ioGPIO_8;
	interface Inout#(Bit#(1)) ioGPIO_9;
	interface Inout#(Bit#(1)) ioGPIO_10;
	interface Inout#(Bit#(1)) ioGPIO_11;
	interface Inout#(Bit#(1)) ioGPIO_12;
	interface Inout#(Bit#(1)) ioGPIO_13;
	interface Inout#(Bit#(1)) ioGPIO_14;
	interface Inout#(Bit#(1)) ioGPIO_15;
	interface Inout#(Bit#(1)) ioI2C1_SCL;
	interface Inout#(Bit#(1)) ioI2C1_SDA;
	interface Inout#(Bit#(1)) ioQSPI0_IO0;
	interface Inout#(Bit#(1)) ioQSPI0_IO1;
	interface Inout#(Bit#(1)) ioQSPI0_IO2;
	interface Inout#(Bit#(1)) ioQSPI0_IO3;
	interface Inout#(Bit#(1)) ioI2C0_SDA;
	interface Inout#(Bit#(1)) ioI2C0_SCL;
	interface Inout#(Bit#(1)) ioSDRAM_D0;
	interface Inout#(Bit#(1)) ioSDRAM_D1;
	interface Inout#(Bit#(1)) ioSDRAM_D2;
	interface Inout#(Bit#(1)) ioSDRAM_D3;
	interface Inout#(Bit#(1)) ioSDRAM_D4;
	interface Inout#(Bit#(1)) ioSDRAM_D5;
	interface Inout#(Bit#(1)) ioSDRAM_D6;
	interface Inout#(Bit#(1)) ioSDRAM_D7;
	interface Inout#(Bit#(1)) ioSDRAM_D8;
	interface Inout#(Bit#(1)) ioSDRAM_D9;
	interface Inout#(Bit#(1)) ioSDRAM_D10;
	interface Inout#(Bit#(1)) ioSDRAM_D11;
	interface Inout#(Bit#(1)) ioSDRAM_D12;
	interface Inout#(Bit#(1)) ioSDRAM_D13;
	interface Inout#(Bit#(1)) ioSDRAM_D14;
	interface Inout#(Bit#(1)) ioSDRAM_D15;
	interface Inout#(Bit#(1)) ioSDRAM_D16;
	interface Inout#(Bit#(1)) ioSDRAM_D17;
	interface Inout#(Bit#(1)) ioSDRAM_D18;
	interface Inout#(Bit#(1)) ioSDRAM_D19;
	interface Inout#(Bit#(1)) ioSDRAM_D20;
	interface Inout#(Bit#(1)) ioSDRAM_D21;
	interface Inout#(Bit#(1)) ioSDRAM_D22;
	interface Inout#(Bit#(1)) ioSDRAM_D23;
	interface Inout#(Bit#(1)) ioSDRAM_D24;
	interface Inout#(Bit#(1)) ioSDRAM_D25;
	interface Inout#(Bit#(1)) ioSDRAM_D26;
	interface Inout#(Bit#(1)) ioSDRAM_D27;
	interface Inout#(Bit#(1)) ioSDRAM_D28;
	interface Inout#(Bit#(1)) ioSDRAM_D29;
	interface Inout#(Bit#(1)) ioSDRAM_D30;
	interface Inout#(Bit#(1)) ioSDRAM_D31;
	method Action iSPI0_MISO (Bit#(1) spi0_mosi);
	method Action iUART0_RX (Bit#(1) uart0_rx);
	method Action iTMS (Bit#(1) tms);
	method Action iTDI (Bit#(1) tdi);
	method Action iSPI1_MISO (Bit#(1) spi1_miso);
	method Action iBOOT_MODE0 (Bit#(1) boot_mode0);
	method Action iBOOT_MODE1 (Bit#(1) boot_mode1);
	method Action iTEST_MODE (Bit#(1) test_mode);
	method Bit#(1) oSPI0_NCS ();
	method Bit#(1) oSPI0_CLK ();
	method Bit#(1) oSPI0_MOSI ();
	method Bit#(1) oQSPI0_CLK ();
	method Bit#(1) oQSPI0_NCS ();
	method Bit#(1) oUART0_TX ();
	method Bit#(1) oTDO ();
	method Bit#(1) oSDRAM_A0 ();
	method Bit#(1) oSDRAM_A1 ();
	method Bit#(1) oSDRAM_A2 ();
	method Bit#(1) oSDRAM_A3 ();
	method Bit#(1) oSDRAM_A4 ();
	method Bit#(1) oSDRAM_A5 ();
	method Bit#(1) oSDRAM_A6 ();
	method Bit#(1) oSDRAM_A7 ();
	method Bit#(1) oSDRAM_A8 ();
	method Bit#(1) oSDRAM_A9 ();
	method Bit#(1) oSDRAM_A10 ();
	method Bit#(1) oSDRAM_A11 ();
	method Bit#(1) oSDRAM_A12 ();
	method Bit#(1) oSDRAM_DQ0 ();
	method Bit#(1) oSDRAM_DQ1 ();
	method Bit#(1) oSDRAM_DQ2 ();
	method Bit#(1) oSDRAM_DQ3 ();
	method Bit#(1) oSDRAM_BA0 ();
	method Bit#(1) oSDRAM_BA1 ();
	method Bit#(1) oSDRAM_CS ();
	method Bit#(1) oSDRAM_RAS ();
	method Bit#(1) oSDRAM_CAS ();
	method Bit#(1) oSDRAM_WE ();
	method Bit#(1) oSDRAM_CLK ();
	method Bit#(1) oSDRAM_CKE ();
	method Bit#(1) oSPI1_NCS ();
	method Bit#(1) oSPI1_CLK ();
	method Bit#(1) oSPI1_MOSI ();
endinterface

import "BVI" aardonyx_wrapper =
module mkaardonyx_wrapper#(Clock iTCK,Reset iTRST)  (Ifc_aardonyx_wrapper);

	default_clock clk_CLK;
	default_reset rst_RESET;

	input_clock clk_CLK (CLK)  <- exposeCurrentClock;
//	input_clock clk_TCK (TCK)  <- tck_CLK;
	input_reset rst_RESET (RESET) clocked_by(clk_CLK)  <- exposeCurrentReset;
	//input_reset rst_TRST (TRST) clocked_by(clk_TCK)  <-trst_RST;

  	ifc_inout ioGPIO_0   (GPIO_0);
	ifc_inout ioGPIO_1   (GPIO_1);       
	ifc_inout ioGPIO_2   (GPIO_2);
	ifc_inout ioGPIO_3   (GPIO_3);
	ifc_inout ioGPIO_4   (GPIO_4);
	ifc_inout ioGPIO_5   (GPIO_5);
	ifc_inout ioGPIO_6   (GPIO_6);
	ifc_inout ioGPIO_7   (GPIO_7);
	ifc_inout ioGPIO_8   (GPIO_8);
	ifc_inout ioGPIO_9   (GPIO_9);
	ifc_inout ioGPIO_10  (GPIO_10);
	ifc_inout ioGPIO_11  (GPIO_11);
	ifc_inout ioGPIO_12  (GPIO_12);
	ifc_inout ioGPIO_13  (GPIO_13);
	ifc_inout ioGPIO_14  (GPIO_14);
	ifc_inout ioGPIO_15  (GPIO_15);
	ifc_inout ioI2C1_SCL (I2C1_SCL);
	ifc_inout ioI2C1_SDA (I2C1_SDA);
	ifc_inout ioQSPI0_IO0(QSPI0_IO0);
	ifc_inout ioQSPI0_IO1(QSPI0_IO1);
	ifc_inout ioQSPI0_IO2(QSPI0_IO2);
	ifc_inout ioQSPI0_IO3(QSPI0_IO3);
	ifc_inout ioI2C0_SDA (I2C0_SDA);
	ifc_inout ioI2C0_SCL (I2C0_SCL);
	ifc_inout ioSDRAM_D0 (SDRAM_D0);
	ifc_inout ioSDRAM_D1 (SDRAM_D1);
	ifc_inout ioSDRAM_D2 (SDRAM_D2);
	ifc_inout ioSDRAM_D3 (SDRAM_D3);
	ifc_inout ioSDRAM_D4 (SDRAM_D4);
	ifc_inout ioSDRAM_D5 (SDRAM_D5);
	ifc_inout ioSDRAM_D6 (SDRAM_D6);
	ifc_inout ioSDRAM_D7 (SDRAM_D7);
	ifc_inout ioSDRAM_D8 (SDRAM_D8);
	ifc_inout ioSDRAM_D9 (SDRAM_D9);
	ifc_inout ioSDRAM_D10(SDRAM_D1);
	ifc_inout ioSDRAM_D11(SDRAM_D1);
	ifc_inout ioSDRAM_D12(SDRAM_D1);
	ifc_inout ioSDRAM_D13(SDRAM_D1);
	ifc_inout ioSDRAM_D14(SDRAM_D1);
	ifc_inout ioSDRAM_D15(SDRAM_D1);
	ifc_inout ioSDRAM_D16(SDRAM_D1);
	ifc_inout ioSDRAM_D17(SDRAM_D1);
	ifc_inout ioSDRAM_D18(SDRAM_D1);
	ifc_inout ioSDRAM_D19(SDRAM_D1);
	ifc_inout ioSDRAM_D20(SDRAM_D2);
	ifc_inout ioSDRAM_D21(SDRAM_D2);
	ifc_inout ioSDRAM_D22(SDRAM_D2);
	ifc_inout ioSDRAM_D23(SDRAM_D2);
	ifc_inout ioSDRAM_D24(SDRAM_D2);
	ifc_inout ioSDRAM_D25(SDRAM_D2);
	ifc_inout ioSDRAM_D26(SDRAM_D2);
	ifc_inout ioSDRAM_D27(SDRAM_D2);
	ifc_inout ioSDRAM_D28(SDRAM_D2);
	ifc_inout ioSDRAM_D29(SDRAM_D2);
	ifc_inout ioSDRAM_D30(SDRAM_D3);
	ifc_inout ioSDRAM_D31(SDRAM_D3);
  

	method iSPI0_MISO (SPI0_MISO)
		 enable((*inhigh*)SPI0_MISO_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iUART0_RX (UART0_RX)
		 enable((*inhigh*)UART0_RX_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iTMS (TMS)
		 enable((*inhigh*)MS_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iTDI (TDI)
		 enable((*inhigh*)TDI_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iSPI1_MISO (SPI1_MISO)
		 enable((*inhigh*)SPI1_MISO_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iBOOT_MODE0 (BOOT_MODE0)
		 enable((*inhigh*)BOOT_MODE0_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iBOOT_MODE1 (BOOT_MODE1)
		 enable((*inhigh*)BOOT_MODE1_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method iTEST_MODE (TEST_MODE)
		 enable((*inhigh*)TEST_MODE_enable) clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI0_NCS oSPI0_NCS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI0_CLK oSPI0_CLK ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI0_MOSI oSPI0_MOSI ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method QSPI0_CLK oQSPI0_CLK ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method QSPI0_NCS oQSPI0_NCS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method UART0_TX oUART0_TX ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method TDO oTDO ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A0 oSDRAM_A0 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A1 oSDRAM_A1 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A2 oSDRAM_A2 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A3 oSDRAM_A3 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A4 oSDRAM_A4 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A5 oSDRAM_A5 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A6 oSDRAM_A6 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A7 oSDRAM_A7 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A8 oSDRAM_A8 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A9 oSDRAM_A9 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A10 oSDRAM_A10 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A11 oSDRAM_A11 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_A12 oSDRAM_A12 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_DQ0 oSDRAM_DQ0 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_DQ1 oSDRAM_DQ1 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_DQ2 oSDRAM_DQ2 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_DQ3 oSDRAM_DQ3 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_BA0 oSDRAM_BA0 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_BA1 oSDRAM_BA1 ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_CS oSDRAM_CS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_RAS oSDRAM_RAS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_CAS oSDRAM_CAS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_WE oSDRAM_WE ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_CLK oSDRAM_CLK ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SDRAM_CKE oSDRAM_CKE ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI1_NCS oSPI1_NCS ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI1_CLK oSPI1_CLK ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);
	method SPI1_MOSI oSPI1_MOSI ()
		 clocked_by(clk_CLK) reset_by(rst_RESET);

	schedule iSPI0_MISO C iSPI0_MISO;
	schedule iSPI0_MISO CF iUART0_RX;
	schedule iSPI0_MISO CF iTMS;
	schedule iSPI0_MISO CF iTDI;
	schedule iSPI0_MISO CF iSPI1_MISO;
	schedule iSPI0_MISO CF iBOOT_MODE0;
	schedule iSPI0_MISO CF iBOOT_MODE1;
	schedule iSPI0_MISO CF iTEST_MODE;
	schedule oSPI0_NCS SB iSPI0_MISO;
	schedule oSPI0_CLK SB iSPI0_MISO;
	schedule oSPI0_MOSI SB iSPI0_MISO;
	schedule oQSPI0_CLK SB iSPI0_MISO;
	schedule oQSPI0_NCS SB iSPI0_MISO;
	schedule oUART0_TX SB iSPI0_MISO;
	schedule oTDO SB iSPI0_MISO;
	schedule oSDRAM_A0 SB iSPI0_MISO;
	schedule oSDRAM_A1 SB iSPI0_MISO;
	schedule oSDRAM_A2 SB iSPI0_MISO;
	schedule oSDRAM_A3 SB iSPI0_MISO;
	schedule oSDRAM_A4 SB iSPI0_MISO;
	schedule oSDRAM_A5 SB iSPI0_MISO;
	schedule oSDRAM_A6 SB iSPI0_MISO;
	schedule oSDRAM_A7 SB iSPI0_MISO;
	schedule oSDRAM_A8 SB iSPI0_MISO;
	schedule oSDRAM_A9 SB iSPI0_MISO;
	schedule oSDRAM_A10 SB iSPI0_MISO;
	schedule oSDRAM_A11 SB iSPI0_MISO;
	schedule oSDRAM_A12 SB iSPI0_MISO;
	schedule oSDRAM_DQ0 SB iSPI0_MISO;
	schedule oSDRAM_DQ1 SB iSPI0_MISO;
	schedule oSDRAM_DQ2 SB iSPI0_MISO;
	schedule oSDRAM_DQ3 SB iSPI0_MISO;
	schedule oSDRAM_BA0 SB iSPI0_MISO;
	schedule oSDRAM_BA1 SB iSPI0_MISO;
	schedule oSDRAM_CS SB iSPI0_MISO;
	schedule oSDRAM_RAS SB iSPI0_MISO;
	schedule oSDRAM_CAS SB iSPI0_MISO;
	schedule oSDRAM_WE SB iSPI0_MISO;
	schedule oSDRAM_CLK SB iSPI0_MISO;
	schedule oSDRAM_CKE SB iSPI0_MISO;
	schedule oSPI1_NCS SB iSPI0_MISO;
	schedule oSPI1_CLK SB iSPI0_MISO;
	schedule oSPI1_MOSI SB iSPI0_MISO;
	schedule iUART0_RX C iUART0_RX;
	schedule iUART0_RX CF iTMS;
	schedule iUART0_RX CF iTDI;
	schedule iUART0_RX CF iSPI1_MISO;
	schedule iUART0_RX CF iBOOT_MODE0;
	schedule iUART0_RX CF iBOOT_MODE1;
	schedule iUART0_RX CF iTEST_MODE;
	schedule oSPI0_NCS SB iUART0_RX;
	schedule oSPI0_CLK SB iUART0_RX;
	schedule oSPI0_MOSI SB iUART0_RX;
	schedule oQSPI0_CLK SB iUART0_RX;
	schedule oQSPI0_NCS SB iUART0_RX;
	schedule oUART0_TX SB iUART0_RX;
	schedule oTDO SB iUART0_RX;
	schedule oSDRAM_A0 SB iUART0_RX;
	schedule oSDRAM_A1 SB iUART0_RX;
	schedule oSDRAM_A2 SB iUART0_RX;
	schedule oSDRAM_A3 SB iUART0_RX;
	schedule oSDRAM_A4 SB iUART0_RX;
	schedule oSDRAM_A5 SB iUART0_RX;
	schedule oSDRAM_A6 SB iUART0_RX;
	schedule oSDRAM_A7 SB iUART0_RX;
	schedule oSDRAM_A8 SB iUART0_RX;
	schedule oSDRAM_A9 SB iUART0_RX;
	schedule oSDRAM_A10 SB iUART0_RX;
	schedule oSDRAM_A11 SB iUART0_RX;
	schedule oSDRAM_A12 SB iUART0_RX;
	schedule oSDRAM_DQ0 SB iUART0_RX;
	schedule oSDRAM_DQ1 SB iUART0_RX;
	schedule oSDRAM_DQ2 SB iUART0_RX;
	schedule oSDRAM_DQ3 SB iUART0_RX;
	schedule oSDRAM_BA0 SB iUART0_RX;
	schedule oSDRAM_BA1 SB iUART0_RX;
	schedule oSDRAM_CS SB iUART0_RX;
	schedule oSDRAM_RAS SB iUART0_RX;
	schedule oSDRAM_CAS SB iUART0_RX;
	schedule oSDRAM_WE SB iUART0_RX;
	schedule oSDRAM_CLK SB iUART0_RX;
	schedule oSDRAM_CKE SB iUART0_RX;
	schedule oSPI1_NCS SB iUART0_RX;
	schedule oSPI1_CLK SB iUART0_RX;
	schedule oSPI1_MOSI SB iUART0_RX;
	schedule iTMS C iTMS;
	schedule iTMS CF iTDI;
	schedule iTMS CF iSPI1_MISO;
	schedule iTMS CF iBOOT_MODE0;
	schedule iTMS CF iBOOT_MODE1;
	schedule iTMS CF iTEST_MODE;
	schedule oSPI0_NCS SB iTMS;
	schedule oSPI0_CLK SB iTMS;
	schedule oSPI0_MOSI SB iTMS;
	schedule oQSPI0_CLK SB iTMS;
	schedule oQSPI0_NCS SB iTMS;
	schedule oUART0_TX SB iTMS;
	schedule oTDO SB iTMS;
	schedule oSDRAM_A0 SB iTMS;
	schedule oSDRAM_A1 SB iTMS;
	schedule oSDRAM_A2 SB iTMS;
	schedule oSDRAM_A3 SB iTMS;
	schedule oSDRAM_A4 SB iTMS;
	schedule oSDRAM_A5 SB iTMS;
	schedule oSDRAM_A6 SB iTMS;
	schedule oSDRAM_A7 SB iTMS;
	schedule oSDRAM_A8 SB iTMS;
	schedule oSDRAM_A9 SB iTMS;
	schedule oSDRAM_A10 SB iTMS;
	schedule oSDRAM_A11 SB iTMS;
	schedule oSDRAM_A12 SB iTMS;
	schedule oSDRAM_DQ0 SB iTMS;
	schedule oSDRAM_DQ1 SB iTMS;
	schedule oSDRAM_DQ2 SB iTMS;
	schedule oSDRAM_DQ3 SB iTMS;
	schedule oSDRAM_BA0 SB iTMS;
	schedule oSDRAM_BA1 SB iTMS;
	schedule oSDRAM_CS SB iTMS;
	schedule oSDRAM_RAS SB iTMS;
	schedule oSDRAM_CAS SB iTMS;
	schedule oSDRAM_WE SB iTMS;
	schedule oSDRAM_CLK SB iTMS;
	schedule oSDRAM_CKE SB iTMS;
	schedule oSPI1_NCS SB iTMS;
	schedule oSPI1_CLK SB iTMS;
	schedule oSPI1_MOSI SB iTMS;
	schedule iTDI C iTDI;
	schedule iTDI CF iSPI1_MISO;
	schedule iTDI CF iBOOT_MODE0;
	schedule iTDI CF iBOOT_MODE1;
	schedule iTDI CF iTEST_MODE;
	schedule oSPI0_NCS SB iTDI;
	schedule oSPI0_CLK SB iTDI;
	schedule oSPI0_MOSI SB iTDI;
	schedule oQSPI0_CLK SB iTDI;
	schedule oQSPI0_NCS SB iTDI;
	schedule oUART0_TX SB iTDI;
	schedule oTDO SB iTDI;
	schedule oSDRAM_A0 SB iTDI;
	schedule oSDRAM_A1 SB iTDI;
	schedule oSDRAM_A2 SB iTDI;
	schedule oSDRAM_A3 SB iTDI;
	schedule oSDRAM_A4 SB iTDI;
	schedule oSDRAM_A5 SB iTDI;
	schedule oSDRAM_A6 SB iTDI;
	schedule oSDRAM_A7 SB iTDI;
	schedule oSDRAM_A8 SB iTDI;
	schedule oSDRAM_A9 SB iTDI;
	schedule oSDRAM_A10 SB iTDI;
	schedule oSDRAM_A11 SB iTDI;
	schedule oSDRAM_A12 SB iTDI;
	schedule oSDRAM_DQ0 SB iTDI;
	schedule oSDRAM_DQ1 SB iTDI;
	schedule oSDRAM_DQ2 SB iTDI;
	schedule oSDRAM_DQ3 SB iTDI;
	schedule oSDRAM_BA0 SB iTDI;
	schedule oSDRAM_BA1 SB iTDI;
	schedule oSDRAM_CS SB iTDI;
	schedule oSDRAM_RAS SB iTDI;
	schedule oSDRAM_CAS SB iTDI;
	schedule oSDRAM_WE SB iTDI;
	schedule oSDRAM_CLK SB iTDI;
	schedule oSDRAM_CKE SB iTDI;
	schedule oSPI1_NCS SB iTDI;
	schedule oSPI1_CLK SB iTDI;
	schedule oSPI1_MOSI SB iTDI;
	schedule iSPI1_MISO C iSPI1_MISO;
	schedule iSPI1_MISO CF iBOOT_MODE0;
	schedule iSPI1_MISO CF iBOOT_MODE1;
	schedule iSPI1_MISO CF iTEST_MODE;
	schedule oSPI0_NCS SB iSPI1_MISO;
	schedule oSPI0_CLK SB iSPI1_MISO;
	schedule oSPI0_MOSI SB iSPI1_MISO;
	schedule oQSPI0_CLK SB iSPI1_MISO;
	schedule oQSPI0_NCS SB iSPI1_MISO;
	schedule oUART0_TX SB iSPI1_MISO;
	schedule oTDO SB iSPI1_MISO;
	schedule oSDRAM_A0 SB iSPI1_MISO;
	schedule oSDRAM_A1 SB iSPI1_MISO;
	schedule oSDRAM_A2 SB iSPI1_MISO;
	schedule oSDRAM_A3 SB iSPI1_MISO;
	schedule oSDRAM_A4 SB iSPI1_MISO;
	schedule oSDRAM_A5 SB iSPI1_MISO;
	schedule oSDRAM_A6 SB iSPI1_MISO;
	schedule oSDRAM_A7 SB iSPI1_MISO;
	schedule oSDRAM_A8 SB iSPI1_MISO;
	schedule oSDRAM_A9 SB iSPI1_MISO;
	schedule oSDRAM_A10 SB iSPI1_MISO;
	schedule oSDRAM_A11 SB iSPI1_MISO;
	schedule oSDRAM_A12 SB iSPI1_MISO;
	schedule oSDRAM_DQ0 SB iSPI1_MISO;
	schedule oSDRAM_DQ1 SB iSPI1_MISO;
	schedule oSDRAM_DQ2 SB iSPI1_MISO;
	schedule oSDRAM_DQ3 SB iSPI1_MISO;
	schedule oSDRAM_BA0 SB iSPI1_MISO;
	schedule oSDRAM_BA1 SB iSPI1_MISO;
	schedule oSDRAM_CS SB iSPI1_MISO;
	schedule oSDRAM_RAS SB iSPI1_MISO;
	schedule oSDRAM_CAS SB iSPI1_MISO;
	schedule oSDRAM_WE SB iSPI1_MISO;
	schedule oSDRAM_CLK SB iSPI1_MISO;
	schedule oSDRAM_CKE SB iSPI1_MISO;
	schedule oSPI1_NCS SB iSPI1_MISO;
	schedule oSPI1_CLK SB iSPI1_MISO;
	schedule oSPI1_MOSI SB iSPI1_MISO;
	schedule iBOOT_MODE0 C iBOOT_MODE0;
	schedule iBOOT_MODE0 CF iBOOT_MODE1;
	schedule iBOOT_MODE0 CF iTEST_MODE;
	schedule oSPI0_NCS SB iBOOT_MODE0;
	schedule oSPI0_CLK SB iBOOT_MODE0;
	schedule oSPI0_MOSI SB iBOOT_MODE0;
	schedule oQSPI0_CLK SB iBOOT_MODE0;
	schedule oQSPI0_NCS SB iBOOT_MODE0;
	schedule oUART0_TX SB iBOOT_MODE0;
	schedule oTDO SB iBOOT_MODE0;
	schedule oSDRAM_A0 SB iBOOT_MODE0;
	schedule oSDRAM_A1 SB iBOOT_MODE0;
	schedule oSDRAM_A2 SB iBOOT_MODE0;
	schedule oSDRAM_A3 SB iBOOT_MODE0;
	schedule oSDRAM_A4 SB iBOOT_MODE0;
	schedule oSDRAM_A5 SB iBOOT_MODE0;
	schedule oSDRAM_A6 SB iBOOT_MODE0;
	schedule oSDRAM_A7 SB iBOOT_MODE0;
	schedule oSDRAM_A8 SB iBOOT_MODE0;
	schedule oSDRAM_A9 SB iBOOT_MODE0;
	schedule oSDRAM_A10 SB iBOOT_MODE0;
	schedule oSDRAM_A11 SB iBOOT_MODE0;
	schedule oSDRAM_A12 SB iBOOT_MODE0;
	schedule oSDRAM_DQ0 SB iBOOT_MODE0;
	schedule oSDRAM_DQ1 SB iBOOT_MODE0;
	schedule oSDRAM_DQ2 SB iBOOT_MODE0;
	schedule oSDRAM_DQ3 SB iBOOT_MODE0;
	schedule oSDRAM_BA0 SB iBOOT_MODE0;
	schedule oSDRAM_BA1 SB iBOOT_MODE0;
	schedule oSDRAM_CS SB iBOOT_MODE0;
	schedule oSDRAM_RAS SB iBOOT_MODE0;
	schedule oSDRAM_CAS SB iBOOT_MODE0;
	schedule oSDRAM_WE SB iBOOT_MODE0;
	schedule oSDRAM_CLK SB iBOOT_MODE0;
	schedule oSDRAM_CKE SB iBOOT_MODE0;
	schedule oSPI1_NCS SB iBOOT_MODE0;
	schedule oSPI1_CLK SB iBOOT_MODE0;
	schedule oSPI1_MOSI SB iBOOT_MODE0;
	schedule iBOOT_MODE1 C iBOOT_MODE1;
	schedule iBOOT_MODE1 CF iTEST_MODE;
	schedule oSPI0_NCS SB iBOOT_MODE1;
	schedule oSPI0_CLK SB iBOOT_MODE1;
	schedule oSPI0_MOSI SB iBOOT_MODE1;
	schedule oQSPI0_CLK SB iBOOT_MODE1;
	schedule oQSPI0_NCS SB iBOOT_MODE1;
	schedule oUART0_TX SB iBOOT_MODE1;
	schedule oTDO SB iBOOT_MODE1;
	schedule oSDRAM_A0 SB iBOOT_MODE1;
	schedule oSDRAM_A1 SB iBOOT_MODE1;
	schedule oSDRAM_A2 SB iBOOT_MODE1;
	schedule oSDRAM_A3 SB iBOOT_MODE1;
	schedule oSDRAM_A4 SB iBOOT_MODE1;
	schedule oSDRAM_A5 SB iBOOT_MODE1;
	schedule oSDRAM_A6 SB iBOOT_MODE1;
	schedule oSDRAM_A7 SB iBOOT_MODE1;
	schedule oSDRAM_A8 SB iBOOT_MODE1;
	schedule oSDRAM_A9 SB iBOOT_MODE1;
	schedule oSDRAM_A10 SB iBOOT_MODE1;
	schedule oSDRAM_A11 SB iBOOT_MODE1;
	schedule oSDRAM_A12 SB iBOOT_MODE1;
	schedule oSDRAM_DQ0 SB iBOOT_MODE1;
	schedule oSDRAM_DQ1 SB iBOOT_MODE1;
	schedule oSDRAM_DQ2 SB iBOOT_MODE1;
	schedule oSDRAM_DQ3 SB iBOOT_MODE1;
	schedule oSDRAM_BA0 SB iBOOT_MODE1;
	schedule oSDRAM_BA1 SB iBOOT_MODE1;
	schedule oSDRAM_CS SB iBOOT_MODE1;
	schedule oSDRAM_RAS SB iBOOT_MODE1;
	schedule oSDRAM_CAS SB iBOOT_MODE1;
	schedule oSDRAM_WE SB iBOOT_MODE1;
	schedule oSDRAM_CLK SB iBOOT_MODE1;
	schedule oSDRAM_CKE SB iBOOT_MODE1;
	schedule oSPI1_NCS SB iBOOT_MODE1;
	schedule oSPI1_CLK SB iBOOT_MODE1;
	schedule oSPI1_MOSI SB iBOOT_MODE1;
	schedule iTEST_MODE C iTEST_MODE;
	schedule oSPI0_NCS SB iTEST_MODE;
	schedule oSPI0_CLK SB iTEST_MODE;
	schedule oSPI0_MOSI SB iTEST_MODE;
	schedule oQSPI0_CLK SB iTEST_MODE;
	schedule oQSPI0_NCS SB iTEST_MODE;
	schedule oUART0_TX SB iTEST_MODE;
	schedule oTDO SB iTEST_MODE;
	schedule oSDRAM_A0 SB iTEST_MODE;
	schedule oSDRAM_A1 SB iTEST_MODE;
	schedule oSDRAM_A2 SB iTEST_MODE;
	schedule oSDRAM_A3 SB iTEST_MODE;
	schedule oSDRAM_A4 SB iTEST_MODE;
	schedule oSDRAM_A5 SB iTEST_MODE;
	schedule oSDRAM_A6 SB iTEST_MODE;
	schedule oSDRAM_A7 SB iTEST_MODE;
	schedule oSDRAM_A8 SB iTEST_MODE;
	schedule oSDRAM_A9 SB iTEST_MODE;
	schedule oSDRAM_A10 SB iTEST_MODE;
	schedule oSDRAM_A11 SB iTEST_MODE;
	schedule oSDRAM_A12 SB iTEST_MODE;
	schedule oSDRAM_DQ0 SB iTEST_MODE;
	schedule oSDRAM_DQ1 SB iTEST_MODE;
	schedule oSDRAM_DQ2 SB iTEST_MODE;
	schedule oSDRAM_DQ3 SB iTEST_MODE;
	schedule oSDRAM_BA0 SB iTEST_MODE;
	schedule oSDRAM_BA1 SB iTEST_MODE;
	schedule oSDRAM_CS SB iTEST_MODE;
	schedule oSDRAM_RAS SB iTEST_MODE;
	schedule oSDRAM_CAS SB iTEST_MODE;
	schedule oSDRAM_WE SB iTEST_MODE;
	schedule oSDRAM_CLK SB iTEST_MODE;
	schedule oSDRAM_CKE SB iTEST_MODE;
	schedule oSPI1_NCS SB iTEST_MODE;
	schedule oSPI1_CLK SB iTEST_MODE;
	schedule oSPI1_MOSI SB iTEST_MODE;
	schedule oSPI0_NCS CF oSPI0_NCS;
	schedule oSPI0_NCS CF oSPI0_CLK;
	schedule oSPI0_NCS CF oSPI0_MOSI;
	schedule oSPI0_NCS CF oQSPI0_CLK;
	schedule oSPI0_NCS CF oQSPI0_NCS;
	schedule oSPI0_NCS CF oUART0_TX;
	schedule oSPI0_NCS CF oTDO;
	schedule oSPI0_NCS CF oSDRAM_A0;
	schedule oSPI0_NCS CF oSDRAM_A1;
	schedule oSPI0_NCS CF oSDRAM_A2;
	schedule oSPI0_NCS CF oSDRAM_A3;
	schedule oSPI0_NCS CF oSDRAM_A4;
	schedule oSPI0_NCS CF oSDRAM_A5;
	schedule oSPI0_NCS CF oSDRAM_A6;
	schedule oSPI0_NCS CF oSDRAM_A7;
	schedule oSPI0_NCS CF oSDRAM_A8;
	schedule oSPI0_NCS CF oSDRAM_A9;
	schedule oSPI0_NCS CF oSDRAM_A10;
	schedule oSPI0_NCS CF oSDRAM_A11;
	schedule oSPI0_NCS CF oSDRAM_A12;
	schedule oSPI0_NCS CF oSDRAM_DQ0;
	schedule oSPI0_NCS CF oSDRAM_DQ1;
	schedule oSPI0_NCS CF oSDRAM_DQ2;
	schedule oSPI0_NCS CF oSDRAM_DQ3;
	schedule oSPI0_NCS CF oSDRAM_BA0;
	schedule oSPI0_NCS CF oSDRAM_BA1;
	schedule oSPI0_NCS CF oSDRAM_CS;
	schedule oSPI0_NCS CF oSDRAM_RAS;
	schedule oSPI0_NCS CF oSDRAM_CAS;
	schedule oSPI0_NCS CF oSDRAM_WE;
	schedule oSPI0_NCS CF oSDRAM_CLK;
	schedule oSPI0_NCS CF oSDRAM_CKE;
	schedule oSPI0_NCS CF oSPI1_NCS;
	schedule oSPI0_NCS CF oSPI1_CLK;
	schedule oSPI0_NCS CF oSPI1_MOSI;
	schedule oSPI0_CLK CF oSPI0_CLK;
	schedule oSPI0_CLK CF oSPI0_MOSI;
	schedule oSPI0_CLK CF oQSPI0_CLK;
	schedule oSPI0_CLK CF oQSPI0_NCS;
	schedule oSPI0_CLK CF oUART0_TX;
	schedule oSPI0_CLK CF oTDO;
	schedule oSPI0_CLK CF oSDRAM_A0;
	schedule oSPI0_CLK CF oSDRAM_A1;
	schedule oSPI0_CLK CF oSDRAM_A2;
	schedule oSPI0_CLK CF oSDRAM_A3;
	schedule oSPI0_CLK CF oSDRAM_A4;
	schedule oSPI0_CLK CF oSDRAM_A5;
	schedule oSPI0_CLK CF oSDRAM_A6;
	schedule oSPI0_CLK CF oSDRAM_A7;
	schedule oSPI0_CLK CF oSDRAM_A8;
	schedule oSPI0_CLK CF oSDRAM_A9;
	schedule oSPI0_CLK CF oSDRAM_A10;
	schedule oSPI0_CLK CF oSDRAM_A11;
	schedule oSPI0_CLK CF oSDRAM_A12;
	schedule oSPI0_CLK CF oSDRAM_DQ0;
	schedule oSPI0_CLK CF oSDRAM_DQ1;
	schedule oSPI0_CLK CF oSDRAM_DQ2;
	schedule oSPI0_CLK CF oSDRAM_DQ3;
	schedule oSPI0_CLK CF oSDRAM_BA0;
	schedule oSPI0_CLK CF oSDRAM_BA1;
	schedule oSPI0_CLK CF oSDRAM_CS;
	schedule oSPI0_CLK CF oSDRAM_RAS;
	schedule oSPI0_CLK CF oSDRAM_CAS;
	schedule oSPI0_CLK CF oSDRAM_WE;
	schedule oSPI0_CLK CF oSDRAM_CLK;
	schedule oSPI0_CLK CF oSDRAM_CKE;
	schedule oSPI0_CLK CF oSPI1_NCS;
	schedule oSPI0_CLK CF oSPI1_CLK;
	schedule oSPI0_CLK CF oSPI1_MOSI;
	schedule oSPI0_MOSI CF oSPI0_MOSI;
	schedule oSPI0_MOSI CF oQSPI0_CLK;
	schedule oSPI0_MOSI CF oQSPI0_NCS;
	schedule oSPI0_MOSI CF oUART0_TX;
	schedule oSPI0_MOSI CF oTDO;
	schedule oSPI0_MOSI CF oSDRAM_A0;
	schedule oSPI0_MOSI CF oSDRAM_A1;
	schedule oSPI0_MOSI CF oSDRAM_A2;
	schedule oSPI0_MOSI CF oSDRAM_A3;
	schedule oSPI0_MOSI CF oSDRAM_A4;
	schedule oSPI0_MOSI CF oSDRAM_A5;
	schedule oSPI0_MOSI CF oSDRAM_A6;
	schedule oSPI0_MOSI CF oSDRAM_A7;
	schedule oSPI0_MOSI CF oSDRAM_A8;
	schedule oSPI0_MOSI CF oSDRAM_A9;
	schedule oSPI0_MOSI CF oSDRAM_A10;
	schedule oSPI0_MOSI CF oSDRAM_A11;
	schedule oSPI0_MOSI CF oSDRAM_A12;
	schedule oSPI0_MOSI CF oSDRAM_DQ0;
	schedule oSPI0_MOSI CF oSDRAM_DQ1;
	schedule oSPI0_MOSI CF oSDRAM_DQ2;
	schedule oSPI0_MOSI CF oSDRAM_DQ3;
	schedule oSPI0_MOSI CF oSDRAM_BA0;
	schedule oSPI0_MOSI CF oSDRAM_BA1;
	schedule oSPI0_MOSI CF oSDRAM_CS;
	schedule oSPI0_MOSI CF oSDRAM_RAS;
	schedule oSPI0_MOSI CF oSDRAM_CAS;
	schedule oSPI0_MOSI CF oSDRAM_WE;
	schedule oSPI0_MOSI CF oSDRAM_CLK;
	schedule oSPI0_MOSI CF oSDRAM_CKE;
	schedule oSPI0_MOSI CF oSPI1_NCS;
	schedule oSPI0_MOSI CF oSPI1_CLK;
	schedule oSPI0_MOSI CF oSPI1_MOSI;
	schedule oQSPI0_CLK CF oQSPI0_CLK;
	schedule oQSPI0_CLK CF oQSPI0_NCS;
	schedule oQSPI0_CLK CF oUART0_TX;
	schedule oQSPI0_CLK CF oTDO;
	schedule oQSPI0_CLK CF oSDRAM_A0;
	schedule oQSPI0_CLK CF oSDRAM_A1;
	schedule oQSPI0_CLK CF oSDRAM_A2;
	schedule oQSPI0_CLK CF oSDRAM_A3;
	schedule oQSPI0_CLK CF oSDRAM_A4;
	schedule oQSPI0_CLK CF oSDRAM_A5;
	schedule oQSPI0_CLK CF oSDRAM_A6;
	schedule oQSPI0_CLK CF oSDRAM_A7;
	schedule oQSPI0_CLK CF oSDRAM_A8;
	schedule oQSPI0_CLK CF oSDRAM_A9;
	schedule oQSPI0_CLK CF oSDRAM_A10;
	schedule oQSPI0_CLK CF oSDRAM_A11;
	schedule oQSPI0_CLK CF oSDRAM_A12;
	schedule oQSPI0_CLK CF oSDRAM_DQ0;
	schedule oQSPI0_CLK CF oSDRAM_DQ1;
	schedule oQSPI0_CLK CF oSDRAM_DQ2;
	schedule oQSPI0_CLK CF oSDRAM_DQ3;
	schedule oQSPI0_CLK CF oSDRAM_BA0;
	schedule oQSPI0_CLK CF oSDRAM_BA1;
	schedule oQSPI0_CLK CF oSDRAM_CS;
	schedule oQSPI0_CLK CF oSDRAM_RAS;
	schedule oQSPI0_CLK CF oSDRAM_CAS;
	schedule oQSPI0_CLK CF oSDRAM_WE;
	schedule oQSPI0_CLK CF oSDRAM_CLK;
	schedule oQSPI0_CLK CF oSDRAM_CKE;
	schedule oQSPI0_CLK CF oSPI1_NCS;
	schedule oQSPI0_CLK CF oSPI1_CLK;
	schedule oQSPI0_CLK CF oSPI1_MOSI;
	schedule oQSPI0_NCS CF oQSPI0_NCS;
	schedule oQSPI0_NCS CF oUART0_TX;
	schedule oQSPI0_NCS CF oTDO;
	schedule oQSPI0_NCS CF oSDRAM_A0;
	schedule oQSPI0_NCS CF oSDRAM_A1;
	schedule oQSPI0_NCS CF oSDRAM_A2;
	schedule oQSPI0_NCS CF oSDRAM_A3;
	schedule oQSPI0_NCS CF oSDRAM_A4;
	schedule oQSPI0_NCS CF oSDRAM_A5;
	schedule oQSPI0_NCS CF oSDRAM_A6;
	schedule oQSPI0_NCS CF oSDRAM_A7;
	schedule oQSPI0_NCS CF oSDRAM_A8;
	schedule oQSPI0_NCS CF oSDRAM_A9;
	schedule oQSPI0_NCS CF oSDRAM_A10;
	schedule oQSPI0_NCS CF oSDRAM_A11;
	schedule oQSPI0_NCS CF oSDRAM_A12;
	schedule oQSPI0_NCS CF oSDRAM_DQ0;
	schedule oQSPI0_NCS CF oSDRAM_DQ1;
	schedule oQSPI0_NCS CF oSDRAM_DQ2;
	schedule oQSPI0_NCS CF oSDRAM_DQ3;
	schedule oQSPI0_NCS CF oSDRAM_BA0;
	schedule oQSPI0_NCS CF oSDRAM_BA1;
	schedule oQSPI0_NCS CF oSDRAM_CS;
	schedule oQSPI0_NCS CF oSDRAM_RAS;
	schedule oQSPI0_NCS CF oSDRAM_CAS;
	schedule oQSPI0_NCS CF oSDRAM_WE;
	schedule oQSPI0_NCS CF oSDRAM_CLK;
	schedule oQSPI0_NCS CF oSDRAM_CKE;
	schedule oQSPI0_NCS CF oSPI1_NCS;
	schedule oQSPI0_NCS CF oSPI1_CLK;
	schedule oQSPI0_NCS CF oSPI1_MOSI;
	schedule oUART0_TX CF oUART0_TX;
	schedule oUART0_TX CF oTDO;
	schedule oUART0_TX CF oSDRAM_A0;
	schedule oUART0_TX CF oSDRAM_A1;
	schedule oUART0_TX CF oSDRAM_A2;
	schedule oUART0_TX CF oSDRAM_A3;
	schedule oUART0_TX CF oSDRAM_A4;
	schedule oUART0_TX CF oSDRAM_A5;
	schedule oUART0_TX CF oSDRAM_A6;
	schedule oUART0_TX CF oSDRAM_A7;
	schedule oUART0_TX CF oSDRAM_A8;
	schedule oUART0_TX CF oSDRAM_A9;
	schedule oUART0_TX CF oSDRAM_A10;
	schedule oUART0_TX CF oSDRAM_A11;
	schedule oUART0_TX CF oSDRAM_A12;
	schedule oUART0_TX CF oSDRAM_DQ0;
	schedule oUART0_TX CF oSDRAM_DQ1;
	schedule oUART0_TX CF oSDRAM_DQ2;
	schedule oUART0_TX CF oSDRAM_DQ3;
	schedule oUART0_TX CF oSDRAM_BA0;
	schedule oUART0_TX CF oSDRAM_BA1;
	schedule oUART0_TX CF oSDRAM_CS;
	schedule oUART0_TX CF oSDRAM_RAS;
	schedule oUART0_TX CF oSDRAM_CAS;
	schedule oUART0_TX CF oSDRAM_WE;
	schedule oUART0_TX CF oSDRAM_CLK;
	schedule oUART0_TX CF oSDRAM_CKE;
	schedule oUART0_TX CF oSPI1_NCS;
	schedule oUART0_TX CF oSPI1_CLK;
	schedule oUART0_TX CF oSPI1_MOSI;
	schedule oTDO CF oTDO;
	schedule oTDO CF oSDRAM_A0;
	schedule oTDO CF oSDRAM_A1;
	schedule oTDO CF oSDRAM_A2;
	schedule oTDO CF oSDRAM_A3;
	schedule oTDO CF oSDRAM_A4;
	schedule oTDO CF oSDRAM_A5;
	schedule oTDO CF oSDRAM_A6;
	schedule oTDO CF oSDRAM_A7;
	schedule oTDO CF oSDRAM_A8;
	schedule oTDO CF oSDRAM_A9;
	schedule oTDO CF oSDRAM_A10;
	schedule oTDO CF oSDRAM_A11;
	schedule oTDO CF oSDRAM_A12;
	schedule oTDO CF oSDRAM_DQ0;
	schedule oTDO CF oSDRAM_DQ1;
	schedule oTDO CF oSDRAM_DQ2;
	schedule oTDO CF oSDRAM_DQ3;
	schedule oTDO CF oSDRAM_BA0;
	schedule oTDO CF oSDRAM_BA1;
	schedule oTDO CF oSDRAM_CS;
	schedule oTDO CF oSDRAM_RAS;
	schedule oTDO CF oSDRAM_CAS;
	schedule oTDO CF oSDRAM_WE;
	schedule oTDO CF oSDRAM_CLK;
	schedule oTDO CF oSDRAM_CKE;
	schedule oTDO CF oSPI1_NCS;
	schedule oTDO CF oSPI1_CLK;
	schedule oTDO CF oSPI1_MOSI;
	schedule oSDRAM_A0 CF oSDRAM_A0;
	schedule oSDRAM_A0 CF oSDRAM_A1;
	schedule oSDRAM_A0 CF oSDRAM_A2;
	schedule oSDRAM_A0 CF oSDRAM_A3;
	schedule oSDRAM_A0 CF oSDRAM_A4;
	schedule oSDRAM_A0 CF oSDRAM_A5;
	schedule oSDRAM_A0 CF oSDRAM_A6;
	schedule oSDRAM_A0 CF oSDRAM_A7;
	schedule oSDRAM_A0 CF oSDRAM_A8;
	schedule oSDRAM_A0 CF oSDRAM_A9;
	schedule oSDRAM_A0 CF oSDRAM_A10;
	schedule oSDRAM_A0 CF oSDRAM_A11;
	schedule oSDRAM_A0 CF oSDRAM_A12;
	schedule oSDRAM_A0 CF oSDRAM_DQ0;
	schedule oSDRAM_A0 CF oSDRAM_DQ1;
	schedule oSDRAM_A0 CF oSDRAM_DQ2;
	schedule oSDRAM_A0 CF oSDRAM_DQ3;
	schedule oSDRAM_A0 CF oSDRAM_BA0;
	schedule oSDRAM_A0 CF oSDRAM_BA1;
	schedule oSDRAM_A0 CF oSDRAM_CS;
	schedule oSDRAM_A0 CF oSDRAM_RAS;
	schedule oSDRAM_A0 CF oSDRAM_CAS;
	schedule oSDRAM_A0 CF oSDRAM_WE;
	schedule oSDRAM_A0 CF oSDRAM_CLK;
	schedule oSDRAM_A0 CF oSDRAM_CKE;
	schedule oSDRAM_A0 CF oSPI1_NCS;
	schedule oSDRAM_A0 CF oSPI1_CLK;
	schedule oSDRAM_A0 CF oSPI1_MOSI;
	schedule oSDRAM_A1 CF oSDRAM_A1;
	schedule oSDRAM_A1 CF oSDRAM_A2;
	schedule oSDRAM_A1 CF oSDRAM_A3;
	schedule oSDRAM_A1 CF oSDRAM_A4;
	schedule oSDRAM_A1 CF oSDRAM_A5;
	schedule oSDRAM_A1 CF oSDRAM_A6;
	schedule oSDRAM_A1 CF oSDRAM_A7;
	schedule oSDRAM_A1 CF oSDRAM_A8;
	schedule oSDRAM_A1 CF oSDRAM_A9;
	schedule oSDRAM_A1 CF oSDRAM_A10;
	schedule oSDRAM_A1 CF oSDRAM_A11;
	schedule oSDRAM_A1 CF oSDRAM_A12;
	schedule oSDRAM_A1 CF oSDRAM_DQ0;
	schedule oSDRAM_A1 CF oSDRAM_DQ1;
	schedule oSDRAM_A1 CF oSDRAM_DQ2;
	schedule oSDRAM_A1 CF oSDRAM_DQ3;
	schedule oSDRAM_A1 CF oSDRAM_BA0;
	schedule oSDRAM_A1 CF oSDRAM_BA1;
	schedule oSDRAM_A1 CF oSDRAM_CS;
	schedule oSDRAM_A1 CF oSDRAM_RAS;
	schedule oSDRAM_A1 CF oSDRAM_CAS;
	schedule oSDRAM_A1 CF oSDRAM_WE;
	schedule oSDRAM_A1 CF oSDRAM_CLK;
	schedule oSDRAM_A1 CF oSDRAM_CKE;
	schedule oSDRAM_A1 CF oSPI1_NCS;
	schedule oSDRAM_A1 CF oSPI1_CLK;
	schedule oSDRAM_A1 CF oSPI1_MOSI;
	schedule oSDRAM_A2 CF oSDRAM_A2;
	schedule oSDRAM_A2 CF oSDRAM_A3;
	schedule oSDRAM_A2 CF oSDRAM_A4;
	schedule oSDRAM_A2 CF oSDRAM_A5;
	schedule oSDRAM_A2 CF oSDRAM_A6;
	schedule oSDRAM_A2 CF oSDRAM_A7;
	schedule oSDRAM_A2 CF oSDRAM_A8;
	schedule oSDRAM_A2 CF oSDRAM_A9;
	schedule oSDRAM_A2 CF oSDRAM_A10;
	schedule oSDRAM_A2 CF oSDRAM_A11;
	schedule oSDRAM_A2 CF oSDRAM_A12;
	schedule oSDRAM_A2 CF oSDRAM_DQ0;
	schedule oSDRAM_A2 CF oSDRAM_DQ1;
	schedule oSDRAM_A2 CF oSDRAM_DQ2;
	schedule oSDRAM_A2 CF oSDRAM_DQ3;
	schedule oSDRAM_A2 CF oSDRAM_BA0;
	schedule oSDRAM_A2 CF oSDRAM_BA1;
	schedule oSDRAM_A2 CF oSDRAM_CS;
	schedule oSDRAM_A2 CF oSDRAM_RAS;
	schedule oSDRAM_A2 CF oSDRAM_CAS;
	schedule oSDRAM_A2 CF oSDRAM_WE;
	schedule oSDRAM_A2 CF oSDRAM_CLK;
	schedule oSDRAM_A2 CF oSDRAM_CKE;
	schedule oSDRAM_A2 CF oSPI1_NCS;
	schedule oSDRAM_A2 CF oSPI1_CLK;
	schedule oSDRAM_A2 CF oSPI1_MOSI;
	schedule oSDRAM_A3 CF oSDRAM_A3;
	schedule oSDRAM_A3 CF oSDRAM_A4;
	schedule oSDRAM_A3 CF oSDRAM_A5;
	schedule oSDRAM_A3 CF oSDRAM_A6;
	schedule oSDRAM_A3 CF oSDRAM_A7;
	schedule oSDRAM_A3 CF oSDRAM_A8;
	schedule oSDRAM_A3 CF oSDRAM_A9;
	schedule oSDRAM_A3 CF oSDRAM_A10;
	schedule oSDRAM_A3 CF oSDRAM_A11;
	schedule oSDRAM_A3 CF oSDRAM_A12;
	schedule oSDRAM_A3 CF oSDRAM_DQ0;
	schedule oSDRAM_A3 CF oSDRAM_DQ1;
	schedule oSDRAM_A3 CF oSDRAM_DQ2;
	schedule oSDRAM_A3 CF oSDRAM_DQ3;
	schedule oSDRAM_A3 CF oSDRAM_BA0;
	schedule oSDRAM_A3 CF oSDRAM_BA1;
	schedule oSDRAM_A3 CF oSDRAM_CS;
	schedule oSDRAM_A3 CF oSDRAM_RAS;
	schedule oSDRAM_A3 CF oSDRAM_CAS;
	schedule oSDRAM_A3 CF oSDRAM_WE;
	schedule oSDRAM_A3 CF oSDRAM_CLK;
	schedule oSDRAM_A3 CF oSDRAM_CKE;
	schedule oSDRAM_A3 CF oSPI1_NCS;
	schedule oSDRAM_A3 CF oSPI1_CLK;
	schedule oSDRAM_A3 CF oSPI1_MOSI;
	schedule oSDRAM_A4 CF oSDRAM_A4;
	schedule oSDRAM_A4 CF oSDRAM_A5;
	schedule oSDRAM_A4 CF oSDRAM_A6;
	schedule oSDRAM_A4 CF oSDRAM_A7;
	schedule oSDRAM_A4 CF oSDRAM_A8;
	schedule oSDRAM_A4 CF oSDRAM_A9;
	schedule oSDRAM_A4 CF oSDRAM_A10;
	schedule oSDRAM_A4 CF oSDRAM_A11;
	schedule oSDRAM_A4 CF oSDRAM_A12;
	schedule oSDRAM_A4 CF oSDRAM_DQ0;
	schedule oSDRAM_A4 CF oSDRAM_DQ1;
	schedule oSDRAM_A4 CF oSDRAM_DQ2;
	schedule oSDRAM_A4 CF oSDRAM_DQ3;
	schedule oSDRAM_A4 CF oSDRAM_BA0;
	schedule oSDRAM_A4 CF oSDRAM_BA1;
	schedule oSDRAM_A4 CF oSDRAM_CS;
	schedule oSDRAM_A4 CF oSDRAM_RAS;
	schedule oSDRAM_A4 CF oSDRAM_CAS;
	schedule oSDRAM_A4 CF oSDRAM_WE;
	schedule oSDRAM_A4 CF oSDRAM_CLK;
	schedule oSDRAM_A4 CF oSDRAM_CKE;
	schedule oSDRAM_A4 CF oSPI1_NCS;
	schedule oSDRAM_A4 CF oSPI1_CLK;
	schedule oSDRAM_A4 CF oSPI1_MOSI;
	schedule oSDRAM_A5 CF oSDRAM_A5;
	schedule oSDRAM_A5 CF oSDRAM_A6;
	schedule oSDRAM_A5 CF oSDRAM_A7;
	schedule oSDRAM_A5 CF oSDRAM_A8;
	schedule oSDRAM_A5 CF oSDRAM_A9;
	schedule oSDRAM_A5 CF oSDRAM_A10;
	schedule oSDRAM_A5 CF oSDRAM_A11;
	schedule oSDRAM_A5 CF oSDRAM_A12;
	schedule oSDRAM_A5 CF oSDRAM_DQ0;
	schedule oSDRAM_A5 CF oSDRAM_DQ1;
	schedule oSDRAM_A5 CF oSDRAM_DQ2;
	schedule oSDRAM_A5 CF oSDRAM_DQ3;
	schedule oSDRAM_A5 CF oSDRAM_BA0;
	schedule oSDRAM_A5 CF oSDRAM_BA1;
	schedule oSDRAM_A5 CF oSDRAM_CS;
	schedule oSDRAM_A5 CF oSDRAM_RAS;
	schedule oSDRAM_A5 CF oSDRAM_CAS;
	schedule oSDRAM_A5 CF oSDRAM_WE;
	schedule oSDRAM_A5 CF oSDRAM_CLK;
	schedule oSDRAM_A5 CF oSDRAM_CKE;
	schedule oSDRAM_A5 CF oSPI1_NCS;
	schedule oSDRAM_A5 CF oSPI1_CLK;
	schedule oSDRAM_A5 CF oSPI1_MOSI;
	schedule oSDRAM_A6 CF oSDRAM_A6;
	schedule oSDRAM_A6 CF oSDRAM_A7;
	schedule oSDRAM_A6 CF oSDRAM_A8;
	schedule oSDRAM_A6 CF oSDRAM_A9;
	schedule oSDRAM_A6 CF oSDRAM_A10;
	schedule oSDRAM_A6 CF oSDRAM_A11;
	schedule oSDRAM_A6 CF oSDRAM_A12;
	schedule oSDRAM_A6 CF oSDRAM_DQ0;
	schedule oSDRAM_A6 CF oSDRAM_DQ1;
	schedule oSDRAM_A6 CF oSDRAM_DQ2;
	schedule oSDRAM_A6 CF oSDRAM_DQ3;
	schedule oSDRAM_A6 CF oSDRAM_BA0;
	schedule oSDRAM_A6 CF oSDRAM_BA1;
	schedule oSDRAM_A6 CF oSDRAM_CS;
	schedule oSDRAM_A6 CF oSDRAM_RAS;
	schedule oSDRAM_A6 CF oSDRAM_CAS;
	schedule oSDRAM_A6 CF oSDRAM_WE;
	schedule oSDRAM_A6 CF oSDRAM_CLK;
	schedule oSDRAM_A6 CF oSDRAM_CKE;
	schedule oSDRAM_A6 CF oSPI1_NCS;
	schedule oSDRAM_A6 CF oSPI1_CLK;
	schedule oSDRAM_A6 CF oSPI1_MOSI;
	schedule oSDRAM_A7 CF oSDRAM_A7;
	schedule oSDRAM_A7 CF oSDRAM_A8;
	schedule oSDRAM_A7 CF oSDRAM_A9;
	schedule oSDRAM_A7 CF oSDRAM_A10;
	schedule oSDRAM_A7 CF oSDRAM_A11;
	schedule oSDRAM_A7 CF oSDRAM_A12;
	schedule oSDRAM_A7 CF oSDRAM_DQ0;
	schedule oSDRAM_A7 CF oSDRAM_DQ1;
	schedule oSDRAM_A7 CF oSDRAM_DQ2;
	schedule oSDRAM_A7 CF oSDRAM_DQ3;
	schedule oSDRAM_A7 CF oSDRAM_BA0;
	schedule oSDRAM_A7 CF oSDRAM_BA1;
	schedule oSDRAM_A7 CF oSDRAM_CS;
	schedule oSDRAM_A7 CF oSDRAM_RAS;
	schedule oSDRAM_A7 CF oSDRAM_CAS;
	schedule oSDRAM_A7 CF oSDRAM_WE;
	schedule oSDRAM_A7 CF oSDRAM_CLK;
	schedule oSDRAM_A7 CF oSDRAM_CKE;
	schedule oSDRAM_A7 CF oSPI1_NCS;
	schedule oSDRAM_A7 CF oSPI1_CLK;
	schedule oSDRAM_A7 CF oSPI1_MOSI;
	schedule oSDRAM_A8 CF oSDRAM_A8;
	schedule oSDRAM_A8 CF oSDRAM_A9;
	schedule oSDRAM_A8 CF oSDRAM_A10;
	schedule oSDRAM_A8 CF oSDRAM_A11;
	schedule oSDRAM_A8 CF oSDRAM_A12;
	schedule oSDRAM_A8 CF oSDRAM_DQ0;
	schedule oSDRAM_A8 CF oSDRAM_DQ1;
	schedule oSDRAM_A8 CF oSDRAM_DQ2;
	schedule oSDRAM_A8 CF oSDRAM_DQ3;
	schedule oSDRAM_A8 CF oSDRAM_BA0;
	schedule oSDRAM_A8 CF oSDRAM_BA1;
	schedule oSDRAM_A8 CF oSDRAM_CS;
	schedule oSDRAM_A8 CF oSDRAM_RAS;
	schedule oSDRAM_A8 CF oSDRAM_CAS;
	schedule oSDRAM_A8 CF oSDRAM_WE;
	schedule oSDRAM_A8 CF oSDRAM_CLK;
	schedule oSDRAM_A8 CF oSDRAM_CKE;
	schedule oSDRAM_A8 CF oSPI1_NCS;
	schedule oSDRAM_A8 CF oSPI1_CLK;
	schedule oSDRAM_A8 CF oSPI1_MOSI;
	schedule oSDRAM_A9 CF oSDRAM_A9;
	schedule oSDRAM_A9 CF oSDRAM_A10;
	schedule oSDRAM_A9 CF oSDRAM_A11;
	schedule oSDRAM_A9 CF oSDRAM_A12;
	schedule oSDRAM_A9 CF oSDRAM_DQ0;
	schedule oSDRAM_A9 CF oSDRAM_DQ1;
	schedule oSDRAM_A9 CF oSDRAM_DQ2;
	schedule oSDRAM_A9 CF oSDRAM_DQ3;
	schedule oSDRAM_A9 CF oSDRAM_BA0;
	schedule oSDRAM_A9 CF oSDRAM_BA1;
	schedule oSDRAM_A9 CF oSDRAM_CS;
	schedule oSDRAM_A9 CF oSDRAM_RAS;
	schedule oSDRAM_A9 CF oSDRAM_CAS;
	schedule oSDRAM_A9 CF oSDRAM_WE;
	schedule oSDRAM_A9 CF oSDRAM_CLK;
	schedule oSDRAM_A9 CF oSDRAM_CKE;
	schedule oSDRAM_A9 CF oSPI1_NCS;
	schedule oSDRAM_A9 CF oSPI1_CLK;
	schedule oSDRAM_A9 CF oSPI1_MOSI;
	schedule oSDRAM_A10 CF oSDRAM_A10;
	schedule oSDRAM_A10 CF oSDRAM_A11;
	schedule oSDRAM_A10 CF oSDRAM_A12;
	schedule oSDRAM_A10 CF oSDRAM_DQ0;
	schedule oSDRAM_A10 CF oSDRAM_DQ1;
	schedule oSDRAM_A10 CF oSDRAM_DQ2;
	schedule oSDRAM_A10 CF oSDRAM_DQ3;
	schedule oSDRAM_A10 CF oSDRAM_BA0;
	schedule oSDRAM_A10 CF oSDRAM_BA1;
	schedule oSDRAM_A10 CF oSDRAM_CS;
	schedule oSDRAM_A10 CF oSDRAM_RAS;
	schedule oSDRAM_A10 CF oSDRAM_CAS;
	schedule oSDRAM_A10 CF oSDRAM_WE;
	schedule oSDRAM_A10 CF oSDRAM_CLK;
	schedule oSDRAM_A10 CF oSDRAM_CKE;
	schedule oSDRAM_A10 CF oSPI1_NCS;
	schedule oSDRAM_A10 CF oSPI1_CLK;
	schedule oSDRAM_A10 CF oSPI1_MOSI;
	schedule oSDRAM_A11 CF oSDRAM_A11;
	schedule oSDRAM_A11 CF oSDRAM_A12;
	schedule oSDRAM_A11 CF oSDRAM_DQ0;
	schedule oSDRAM_A11 CF oSDRAM_DQ1;
	schedule oSDRAM_A11 CF oSDRAM_DQ2;
	schedule oSDRAM_A11 CF oSDRAM_DQ3;
	schedule oSDRAM_A11 CF oSDRAM_BA0;
	schedule oSDRAM_A11 CF oSDRAM_BA1;
	schedule oSDRAM_A11 CF oSDRAM_CS;
	schedule oSDRAM_A11 CF oSDRAM_RAS;
	schedule oSDRAM_A11 CF oSDRAM_CAS;
	schedule oSDRAM_A11 CF oSDRAM_WE;
	schedule oSDRAM_A11 CF oSDRAM_CLK;
	schedule oSDRAM_A11 CF oSDRAM_CKE;
	schedule oSDRAM_A11 CF oSPI1_NCS;
	schedule oSDRAM_A11 CF oSPI1_CLK;
	schedule oSDRAM_A11 CF oSPI1_MOSI;
	schedule oSDRAM_A12 CF oSDRAM_A12;
	schedule oSDRAM_A12 CF oSDRAM_DQ0;
	schedule oSDRAM_A12 CF oSDRAM_DQ1;
	schedule oSDRAM_A12 CF oSDRAM_DQ2;
	schedule oSDRAM_A12 CF oSDRAM_DQ3;
	schedule oSDRAM_A12 CF oSDRAM_BA0;
	schedule oSDRAM_A12 CF oSDRAM_BA1;
	schedule oSDRAM_A12 CF oSDRAM_CS;
	schedule oSDRAM_A12 CF oSDRAM_RAS;
	schedule oSDRAM_A12 CF oSDRAM_CAS;
	schedule oSDRAM_A12 CF oSDRAM_WE;
	schedule oSDRAM_A12 CF oSDRAM_CLK;
	schedule oSDRAM_A12 CF oSDRAM_CKE;
	schedule oSDRAM_A12 CF oSPI1_NCS;
	schedule oSDRAM_A12 CF oSPI1_CLK;
	schedule oSDRAM_A12 CF oSPI1_MOSI;
	schedule oSDRAM_DQ0 CF oSDRAM_DQ0;
	schedule oSDRAM_DQ0 CF oSDRAM_DQ1;
	schedule oSDRAM_DQ0 CF oSDRAM_DQ2;
	schedule oSDRAM_DQ0 CF oSDRAM_DQ3;
	schedule oSDRAM_DQ0 CF oSDRAM_BA0;
	schedule oSDRAM_DQ0 CF oSDRAM_BA1;
	schedule oSDRAM_DQ0 CF oSDRAM_CS;
	schedule oSDRAM_DQ0 CF oSDRAM_RAS;
	schedule oSDRAM_DQ0 CF oSDRAM_CAS;
	schedule oSDRAM_DQ0 CF oSDRAM_WE;
	schedule oSDRAM_DQ0 CF oSDRAM_CLK;
	schedule oSDRAM_DQ0 CF oSDRAM_CKE;
	schedule oSDRAM_DQ0 CF oSPI1_NCS;
	schedule oSDRAM_DQ0 CF oSPI1_CLK;
	schedule oSDRAM_DQ0 CF oSPI1_MOSI;
	schedule oSDRAM_DQ1 CF oSDRAM_DQ1;
	schedule oSDRAM_DQ1 CF oSDRAM_DQ2;
	schedule oSDRAM_DQ1 CF oSDRAM_DQ3;
	schedule oSDRAM_DQ1 CF oSDRAM_BA0;
	schedule oSDRAM_DQ1 CF oSDRAM_BA1;
	schedule oSDRAM_DQ1 CF oSDRAM_CS;
	schedule oSDRAM_DQ1 CF oSDRAM_RAS;
	schedule oSDRAM_DQ1 CF oSDRAM_CAS;
	schedule oSDRAM_DQ1 CF oSDRAM_WE;
	schedule oSDRAM_DQ1 CF oSDRAM_CLK;
	schedule oSDRAM_DQ1 CF oSDRAM_CKE;
	schedule oSDRAM_DQ1 CF oSPI1_NCS;
	schedule oSDRAM_DQ1 CF oSPI1_CLK;
	schedule oSDRAM_DQ1 CF oSPI1_MOSI;
	schedule oSDRAM_DQ2 CF oSDRAM_DQ2;
	schedule oSDRAM_DQ2 CF oSDRAM_DQ3;
	schedule oSDRAM_DQ2 CF oSDRAM_BA0;
	schedule oSDRAM_DQ2 CF oSDRAM_BA1;
	schedule oSDRAM_DQ2 CF oSDRAM_CS;
	schedule oSDRAM_DQ2 CF oSDRAM_RAS;
	schedule oSDRAM_DQ2 CF oSDRAM_CAS;
	schedule oSDRAM_DQ2 CF oSDRAM_WE;
	schedule oSDRAM_DQ2 CF oSDRAM_CLK;
	schedule oSDRAM_DQ2 CF oSDRAM_CKE;
	schedule oSDRAM_DQ2 CF oSPI1_NCS;
	schedule oSDRAM_DQ2 CF oSPI1_CLK;
	schedule oSDRAM_DQ2 CF oSPI1_MOSI;
	schedule oSDRAM_DQ3 CF oSDRAM_DQ3;
	schedule oSDRAM_DQ3 CF oSDRAM_BA0;
	schedule oSDRAM_DQ3 CF oSDRAM_BA1;
	schedule oSDRAM_DQ3 CF oSDRAM_CS;
	schedule oSDRAM_DQ3 CF oSDRAM_RAS;
	schedule oSDRAM_DQ3 CF oSDRAM_CAS;
	schedule oSDRAM_DQ3 CF oSDRAM_WE;
	schedule oSDRAM_DQ3 CF oSDRAM_CLK;
	schedule oSDRAM_DQ3 CF oSDRAM_CKE;
	schedule oSDRAM_DQ3 CF oSPI1_NCS;
	schedule oSDRAM_DQ3 CF oSPI1_CLK;
	schedule oSDRAM_DQ3 CF oSPI1_MOSI;
	schedule oSDRAM_BA0 CF oSDRAM_BA0;
	schedule oSDRAM_BA0 CF oSDRAM_BA1;
	schedule oSDRAM_BA0 CF oSDRAM_CS;
	schedule oSDRAM_BA0 CF oSDRAM_RAS;
	schedule oSDRAM_BA0 CF oSDRAM_CAS;
	schedule oSDRAM_BA0 CF oSDRAM_WE;
	schedule oSDRAM_BA0 CF oSDRAM_CLK;
	schedule oSDRAM_BA0 CF oSDRAM_CKE;
	schedule oSDRAM_BA0 CF oSPI1_NCS;
	schedule oSDRAM_BA0 CF oSPI1_CLK;
	schedule oSDRAM_BA0 CF oSPI1_MOSI;
	schedule oSDRAM_BA1 CF oSDRAM_BA1;
	schedule oSDRAM_BA1 CF oSDRAM_CS;
	schedule oSDRAM_BA1 CF oSDRAM_RAS;
	schedule oSDRAM_BA1 CF oSDRAM_CAS;
	schedule oSDRAM_BA1 CF oSDRAM_WE;
	schedule oSDRAM_BA1 CF oSDRAM_CLK;
	schedule oSDRAM_BA1 CF oSDRAM_CKE;
	schedule oSDRAM_BA1 CF oSPI1_NCS;
	schedule oSDRAM_BA1 CF oSPI1_CLK;
	schedule oSDRAM_BA1 CF oSPI1_MOSI;
	schedule oSDRAM_CS CF oSDRAM_CS;
	schedule oSDRAM_CS CF oSDRAM_RAS;
	schedule oSDRAM_CS CF oSDRAM_CAS;
	schedule oSDRAM_CS CF oSDRAM_WE;
	schedule oSDRAM_CS CF oSDRAM_CLK;
	schedule oSDRAM_CS CF oSDRAM_CKE;
	schedule oSDRAM_CS CF oSPI1_NCS;
	schedule oSDRAM_CS CF oSPI1_CLK;
	schedule oSDRAM_CS CF oSPI1_MOSI;
	schedule oSDRAM_RAS CF oSDRAM_RAS;
	schedule oSDRAM_RAS CF oSDRAM_CAS;
	schedule oSDRAM_RAS CF oSDRAM_WE;
	schedule oSDRAM_RAS CF oSDRAM_CLK;
	schedule oSDRAM_RAS CF oSDRAM_CKE;
	schedule oSDRAM_RAS CF oSPI1_NCS;
	schedule oSDRAM_RAS CF oSPI1_CLK;
	schedule oSDRAM_RAS CF oSPI1_MOSI;
	schedule oSDRAM_CAS CF oSDRAM_CAS;
	schedule oSDRAM_CAS CF oSDRAM_WE;
	schedule oSDRAM_CAS CF oSDRAM_CLK;
	schedule oSDRAM_CAS CF oSDRAM_CKE;
	schedule oSDRAM_CAS CF oSPI1_NCS;
	schedule oSDRAM_CAS CF oSPI1_CLK;
	schedule oSDRAM_CAS CF oSPI1_MOSI;
	schedule oSDRAM_WE CF oSDRAM_WE;
	schedule oSDRAM_WE CF oSDRAM_CLK;
	schedule oSDRAM_WE CF oSDRAM_CKE;
	schedule oSDRAM_WE CF oSPI1_NCS;
	schedule oSDRAM_WE CF oSPI1_CLK;
	schedule oSDRAM_WE CF oSPI1_MOSI;
	schedule oSDRAM_CLK CF oSDRAM_CLK;
	schedule oSDRAM_CLK CF oSDRAM_CKE;
	schedule oSDRAM_CLK CF oSPI1_NCS;
	schedule oSDRAM_CLK CF oSPI1_CLK;
	schedule oSDRAM_CLK CF oSPI1_MOSI;
	schedule oSDRAM_CKE CF oSDRAM_CKE;
	schedule oSDRAM_CKE CF oSPI1_NCS;
	schedule oSDRAM_CKE CF oSPI1_CLK;
	schedule oSDRAM_CKE CF oSPI1_MOSI;
	schedule oSPI1_NCS CF oSPI1_NCS;
	schedule oSPI1_NCS CF oSPI1_CLK;
	schedule oSPI1_NCS CF oSPI1_MOSI;
	schedule oSPI1_CLK CF oSPI1_CLK;
	schedule oSPI1_CLK CF oSPI1_MOSI;
	schedule oSPI1_MOSI CF oSPI1_MOSI;
endmodule


